��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}����Q%b<Y�D&�u�"��U���T��ײ2��>���^k�/7�?1�(�c��ߘ�]��|�G��f�:��#tC��o�Rb�v �mD�?�D��L���_�L����\�Q^������*r���`���N�w	*D���y&�f��+K��[y��ڂ�Vs>�+���,>z���/lt�3� P�;��1�-��⫯g*P(�C#<�:z����uP!ߌ��˼�{�&�z(ݲm@��Q��D(
b�r�5�c$e
�9��Ax!P�����M~�-~����U��[��LUP4��R  ���~��X�F�n� )�\�~xy����"�L���om�Q*���T�K/ZT�@�(X!��N��j�㝣�Ĭ�Jn�ru�����&��5|��Հ��qyA��f
�,�;��w�AV��'}�F�b_r��'�Y�a��s���M�.ѳ��b��NmJ0i�,�L�R�b���T�g���#Zm�|foV�v�^U�v��8@8ز�󟾏�{A��Y���4IQm��*b.[P��1��+n$�̇���S~$�}>���8��0�uw���j������x��(���a���<5(N����7W-��L�@�y����L
�T�p r��|���-&�TfH8E^���G�H�8|�0?�+�~c(�"��Y��q s�y�(�������2�#,�Է/�o�po���1�]�����u�)[9{��5.V��ȍ�gj���K�X`��_/�ߏ����89!#1l���=?��nnD6�!��հI#ķ�/T�ʭ��<?�9}�Ƿ���WE�-��mD>�0a���/�w�'Oq��w��`Y�s�J�0o��
�m�᢯��0���6=�[�߹� @�S���Q��G��l*&p�Yy�yB�򊓳q9M38���E�!���<< �sN۪�c�	u�~Rp�,k���%k�&ָ��sE��D�őⴔIꈸV�MT7xB2I�d�HnULkIh��:h
�[ϸ��W�A��S;CM���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc(#`��Gcp��}K��f<�,=K�F~�?|�[_X��ˆk�=�sQ��X�zȣc��- ��Ckӏ�^!�:�_c�~:i��p�7��Xi9�
�ѹaB��Q�//?�s�m/C�N{a�9O!JoE'U�Y�y��
r�)�Y¹w����i��T!R����.�D���J7"H�f�J2�ѬL�1m��+Y#_WӢۉ���2=�l�����뙇�� E�{���_�-h|,���(����>S��ә�����/�4�}n'���a*�x���� ����ޙB!7����ˉ�1�:�Ω�s8�R�	�}����Q%b<Y�D�IY��L�Π��Ǣ&�3ݾw�����$G⃍�����i3<�f�D���X���`��wl��h��"u����i��؞��b9����{oS�2>� zM�Xh�hk�i��i���'n�^0o�h{4N'�Ī���������aIXƕ{�������®�������S���ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3|^�3�]�h}ZJB�����r)4qA��oj��n���k���{7$0~'��Qv�)�o��:�zL͊�q��1�KB|1<\��D?��Ǳ�0|]<w:�>���'hZ���j�Q%��{S'�����E�E)�6����#±�sR�{F;�f��X�����.��7bAg�
d�m�Zu�P�{@���u��7+��ا��,�!�`�(i3!�`�(i3!�`�(i3!�`�(i3� ͷ�	�~�J�_�Ď	��[�!%]���A�����y������i�=]A��O�T=�4e=��-������yMK�o�Y�Q�;�Q+�[Z��=]A��O�T=�4e=��-�*&�[��/���i� �j[�YP����M�g����!�`�(i3v�ј�"��Z鎬�����X���*�V��*J "�,�>E����-��%Mό���.� ���M��2�����Vc�q`<�5W�Օq�]�ŀ!0��Á�j*�tߪ��a#�f�E����F7G#+�Ǘ0z�cUL��Jv(K�V��W��_�ړ8���/��P���w��:
1���Ɣw��/w~���j��3L��'9�*�p9��b�^��\��[|��w��T�mT\-!�`�(i3!�`�(i3!�`�(i3!�`�(i3%m�\�u��I�z�]NW���:j���Բv�+@!�`�(i3!�`�(i3!�`�(i3!�`�(i3D�k���?�8c�	�^�贅����	^�������!�m���d��E����F7G#+��3L��'9�O�^Q��h���LDY�P|�gd#v�5�!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=WlF��8�j�6G���8i�qcU������~�A�qIp��K�ӅKW@IE�U����S8�bM� 2)G��8���/���\Zd�O���&z��&����壃�b��'����R�c�ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3Bq�`c�!1�b[����J�-Kѐ�f�U-I�g_$?��uk0!�`�(i3!�`�(i3!�`�(i3!�`�(i3���y��lDKw�UnM��H��(.�gPbT8�����9��s+"��n�I�7�p�����E��@IE�U��`�-9v��"�����B�K��L!b!��u�4�����7J|et����$!�`�(i3!�`�(i3!�`�(i3!�`�(i3���y��lD���bxA�����|*>i�ܻ��`���&U������J z͝�1y�<.��2-"�,�>E���TD��-�`��8�4P�d�=/;����T�a����]Q�ߣ�b2�{��OJ<�a��d�ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�/[��� ����=6�p}���*_����s5�����D�pc�2�����VcaC����:��I�e�öZr
�0�M�yObFT+V������P.g"}�p�Ԭ����
L'���Xwa�Ĝz�n~�r%ӷ��#�jV�����Sw�l6�P��{�!�`�(i3!�`�(i3!�`�(i3!�`�(i3Wݡ������!�qgGq�% �-;�(��v��%��������P�A������|g�Y�'���Xw�.aX�bAK��U�,��/��K�*� ���j���0z�cUL��Jv(K�V��W��_�ړ8���/��.aX�bAKJ0i�,�L����_����j��<ͧ�:|��b+}y[����C=+f5��pw�b�v�ј�"��Z鎬����Ĺ#{���.aX�bAK����e_��':E����j���0z�cUL���.�1�3�8���/�Յ՝a��h�JE�(����X%���ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�R�����3�����t,G넗]��D�Y��0���R]�K����cg��tӱ1R�m��+�<4��ˌ�ň��h��֑�/6K�R�8�bϣ��'�����N<���d�k��Yu>�G Oag�qod�֓��+��T���jB�Fg�Y씤`��p�܂aQ�l&K[�
C&����k�+ND�A���@�k��V�4���|;��7����Re�.QZ�$ą_�����D�**����W�fYCJd<���FuIL�; � e�m���Ը
�7���f�,,�2���7#[+��z�6̇"�W��@�Aw��1���mr���h''�I�َG����PE��I��'������[��CCLn��S�W#w���	(���B�� ��I�=M�^"4/�������*���I��'�!͙��04nry��cT���D	��U�l>o��|�=���yp�.P��&��c=T7fÃl����4�,�dט�w���rvZ�b��^���B0S�=�א=ͼ�\�vś��X&`�Kb�����=gA���_5p}w>���uS ��������s�0F1��D�I�t�5����`Ko�F)���;4����)\|�^��
�>IÙ=�H���]*����*Tt���#��0u���%��0�P������qθO.�r���$��^��Bcƕrͼ���\����iW5�z�a$��u1#��Z�����XP��ȬvbëdP`����Oh����w�G��^��ه�U�Yyr��$d�I�v�|��lX�.8o�A����5�e`��9̖UB�no�B��+ Hxg`�H�4��`t�A~�@����gG�Q�e��)Z���_j���M"��q����Oއ�?t},�׉é[�=�5x�зq.|KH�"�,�>E���]�!���e��Ƥ����n9�F�,g�ul7����n`5�fK�\w��0]7��"=��<D�n:3MO�`�Wi&����i�#Ѻ'���Xw���,D���`��/s�1��pзq8�Ј'���Xw���,D\X��!��^�T�H���зq8�Ј'���Xw���,D\X��!��!�`�(i3��lJ��튝�b�Bϱ������[��CC��a�(��R�wX��}�
�?���v�)y�Eh�ѮYțx z�Jm]�#�;� ��B�D�F ���~=�L�����3��7s�9���o>��l%i�-}ϼ 8����Ƀ�?PA�g�+C��s7s�9���o��S8�bM� 2)G��8���/����,Dߔ��� �3y��5����'���Xw�j�7��a(􆿳����d/h�5�G�G�����y���Υ�d[g��Q]� _ό���.�}�
�?�������P�]Z������Q]� _ό���.�}�
�?�������P�8�>�}���Q]� _ό���.��7�b�������6}G�?-�D�E����FZ鎬�������*�n�B.W���ۗ$|�N
�`!�`�(i37s�9���o!��w���J*��9W���bv���H˳͠m�xW��-#��k+m�&���w/s�!g#��������WT� �`�o��)��.��!�`�(i3�d�٣���N N�S��E �����VF�˷�!�`�(i3�d�٣���N N�S��E �����VF�˷�BڴQ���n`5�fK�\w��0]7��"=��T��+𦊢~�s��9����+�J���q���U��@����gG�m�n�~�!�G���-���+�J���q���U��˞�Bx�i�p��+�PUѦ�Ƴ��a�W�Z鎬�������*�n�B�E ����*{��[�$�!�`�(i3�d�٣���N N�S�D[��+s�c�~$幙xn����U'�q���U��@����gG�8��y�l�H����I�d�٣��4�5_�o0b!��u��΁M�$���� B�J���]�!����-ዧ�[����n9�������(ݝWu/k��Z鎬��������l��:|m1�_^c���\�X7s�9���o>��l%i�-5�e`��94\%��t�,�Qy*ό���.�aZ��qA�EFmғO�4}�G��зq8�Ј'���Xw���,DFmғO�4}`L����D:зq8�Ј'���Xw���,DFmғO�4}5���u�L���Q]� _�rs�i���`�M�	=̞��>��vbëdP�D�R��	ܷ�4D�P~��#��#��T�\ ���ό�]2�E ����cݵ�Ǡ��0���Y$��d�٣���o��D���/h�5�G�G��2�b=�e���b��n`5�fK��0z�cUL��Jv(K�V��W��_�ړ8���/����,D�d^�-Z?�������(���G
'���Xw�j�7���5�%]���a(􆿳���2����.��g#���7�|�[�A�J�d�٣���N N�S���g#���7�|'!�b9���d�٣���N N�S�	�:-!@xNm���d���Υ�d[g�d�٣���N N�S�	�:-!@xNm���d�=�������d�٣���N N�S��E ����Z���]�}�zM#��m��d�٣��c�A�L'������ڂ�ޕR�wX��}�
�?�Vi� �ZD�o�&��Q]� _�rs�i��s�٭����D�h��T�\ ��i3�|)sՀ/�n�*���e���b��E����FZ鎬�����
!-�n����b��yt��\�Dk���|WLP|��#��ZBi�mR!.<ή�$	�:-!@xN ��\�&ɖ��_j���	�k���	�U���q�
�ep�G;w�b!��u�g�G��0�2 �����ό���.�}�
�?���"���l<o�;)�y�y�����d�٣���o��D���/h�5�G�G�M��L�%�1�@ �~)�d�٣���N N�S���z@�����E��B�1� �-5$�w=����d�.��j�ـ���Qgă�����󼻄��Lv����M1��:O��_�:��K'*|����7�|�[�A�J� 	��^��뒋N�nX�8jUG�*"���6Bj�!�`�(i3!�`�(i3�ٿ�^���u�p��;�����U�-��h��ڥ����Ⱦy:Ɔ�P�oX��Q��eV#GS�܇5*A�u����l0����'{w#/ B!�`�(i3!�`�(i3�����ziT˗=߫����L$�$���8�5�b��+N���ˇmWᅫw�5�O�%E#P}�
�?�i�:`�+P_2�
C�]�!��`��j(&�L��K��I/N#~8"�Z�z��B��������p���?U��zC�4M/�Sн3y��
~i�g����8���b�2�w�����-����/T�=qއ*|�ވQ�:� 	��^�Bg�1�/?~$�}>���w�q����gVdxQ,�<@���ل=����h�)N�'n�쮾�\�i\!�`�(i3!�`�(i3�V.9��L=�q��G8��"[�GVg��x�����{���������EN.<��{��x� I,��̖UB�no�d�;�����6Bj�!�`�(i3!�`�(i3�����z΃/��}�y6�T�@�����L�6�o8:4�g�G��0>߰�e��A�Ҷ����Sl��!�`�(i3!�`�(i3!�`�(i3��'T���+��e�D.7�gqSά�B�����e_�,9�f��������P�꠼*d�m?�#	*]]�iI9�o«IX0F�M��Eg�뚵]k�WM��q|���N�ui����0K�~���`UNP�G�&ց�*�#�vzR5�<���>e�-�����@:[�X)P<�ܓ�Y!�`�(i3@v��e��~$�}>���w�q���_�mS8<�n�ݚ�Н��7����������EN.74/���g!�%=F�=!�`�(i3�����!�`�(i3���g!h!���7�|���޵.�۬gVdxQ,�K��I/��0�|��';��#j�ݚ�Н���+�t2��Lq��QF[��f�\%���}��ݚ�Н��Ra])n#]���\�x8�:
1����0/0`9N1>!XM�#����+1�;�.��1���-����!�`�(i3�D�������{
Bk	䶙%T7u��2�!�`�(i3�k��^�1�K��I/z�
1���;#o�]�ʄ�
%�6W���N�Cٺ��������� h�ҩ�!�`�(i3@��( ���M/*�3�s��m�Eq�e>%����
�:qEp���,��\[��l�,t���H[W?��v[v%���e�D.7�q���f�e�M?��y�!�`�(i3����&��r��졾�g�Y���v�l���"!�`�(i3��w�w:�!�`�(i3����&��r��졾�g�Y�٩�����ݚ�Н�fĉ>99��A0ok��
�:qEp�;�P�t�5��6��UH6"����K˖�s9�O��F����{L,84a��|�&��}Dq�f���Aڬ&W럼�~=�L�����3���'����u��r��!�`�(i3�<@���ل=����h�Wsp[��X��=@'ѥ��Ra])n#���r����;�jmT�#������P�꠼*d�m1F#�֞qduP���2
�M����d9=���u��r��!�`�(i3h5���=�t���_j���Gƻ������Ɇ�5�!�`�(i3��\7�fˁ��7�|���޵.�۬gVdxQ,�K��I/��0�|�_�mS8<�n�ݚ�Н���+�t2��Lq��QF[��f�\%���}��ݚ�Н��Ra])n#]���\�x8�:
1���Ư����z��>!XM�#����+1��*Hx�g���-����!�`�(i3�D�������{
Bk	䶙%�+���q��!�`�(i3�k��^�1�K��I/z�
1���;#o�]�ʄ�
%�6W���N�Cٺ��G��Hb� h�ҩ�!�`�(i3@��( ���M/*�3��{��3���}Dq�f�՝� s�#���k$ !�`�(i3@��( ���M/*�3����3��[<�m��I�!�`�(i3�5ߧE4��!�`�(i3��Ě���ž_�F�(*�O�q�u�PH<!�`�(i3�U�Z^�t� "���
w���NM�������l��T���ӄ`^�Ad0t�;!��Q�����&G!�`�(i3�o�t����w�`L����Y� �K;��t��:!�`�(i31���~!�`�(i3@v��e��֯���,�ۿ���L��:����iW3��O�����%�������&G!�`�(i3�7����������EN.74/������.ݍ|�!�`�(i3�̢k���������P�꠼*d�m1F#�֞qduP���2
�M����'����u��r��!�`�(i3h5���=�t���_j���Gƻ������Ɇ�5�!�`�(i3��\7�fˁ��7�|���޵.�ۃVa�ir�K��I/��0�|��';��#j�ݚ�Н���+�t2��Lq��QF[��f�\%h���UZ���ݚ�Н��Ra])n#]���\�x8�:
1���Ư����z��>!XM�#����+1�;�.��1���-����!�`�(i3�D�������{
B֗M-k��%)z�
3Me!�`�(i3��jVѭ@!�`�(i3�D�������{
Bk	䶙%G�kk�!�`�(i3$f��_Ub�F�S�1 �fĉ>99��j���Gp�ݓ�W���=�����]s���D*j9�O��F����{L,84a��|�&��}Dq�f���Aڬ&W럼�~=�L�����3���'����u��r��!�`�(i3�<@���ل=����h�Wsp[��X��=@'ѥ��Ra])n#���r����;�jmT�#������P�꠼*d�m1F#�֞qduP���2
�M����d9=���u��r��!�`�(i3h5���=�t���_j���Gƻ������Ɇ�5�!�`�(i3��\7�fˁ��7�|���޵.�۬gVdxQ,�K��I/��0�|�_�mS8<�n�ݚ�Н���+�t2��Lq��QF[��f�\%���}��ݚ�Н��Ra])n#]���\�x8�:
1���Ư����z��>!XM�#����+1��*Hx�g���-����!�`�(i3�D�������{
Bk	䶙%�+���q��!�`�(i3�k��^�1�K��I/z�
1���;#o�]�ʄ�
%�6W���N�Cٺ��G��Hb� h�ҩ�!�`�(i3@��( ���M/*�3��{��3���}Dq�f�՝� s�#���k$ !�`�(i3@��( ���M/*�3����3��[<�m��I�!�`�(i3�5ߧE4��!�`�(i3��Ě���ž_�F�(*�O�qe��0�U���>e�D�������{
Bk	䶙%G�kk�!�`�(i3���4)c-�¾L���q9+t�}�;b�-�2��Q������}�	76�&�φ��<�6�U�7˖�ɳ
xM�v.���������,�ǰ����ԫ�`RO���֑I�_D��L��ީ)�G�h�4n�9gl�	�Q
��?��u��"u����:/�)0�/���H�V���羹��K��I/N#~8"�Z�z��B��������p��DO&��N������Px"S�#�d+�_0c �6�_ܸy^�J����p�@OM.Ir���UHf�����_j����d�;��-͍�Ձo��{
B���ͽ�n-=�,�*ːD�f�.��!�`�(i3!�`�(i3��r-��r��졾�g��[��o}���p������6Bj�!�`�(i3!�`�(i3}Y;�jn��|��p���˃�I��x���_��.)<�ʮ�{
BfxQ�-V�N|~�.�u���r����!�`�(i3��7I����4��}�<�"[�GVg��x���_��.)<�ʮ�{
BX{J�[�,uM[x7i��r��졾�g��[��o}���O�!�`�(i3!�`�(i3Lz8�D��<��{��x� I,��̖UB�no �ilچ=���6Bj�!�`�(i3!�`�(i3/��kOT��3�l�=�K����
]�vp����t�T��4c�� n�ƫ�}<��K��I/�x���L�������P����݀e�O��z%�ԬQ���&���贵!�`�(i3!�`�(i3!�`�(i3��F�������p�,���:���~$�}>����k`�Ӊ�'���>;#M�"����!�`�(i3!�`�(i3!�`�(i3�_��>νr�T�g���:�0��7#�z�3��#���n?�#	*]]�iI9�o«IX0F�M��Eg�뚵]k�WM��q!��p4��ui����0K�~���`UNP�G�&ց�*�#�vzR5�<���>e�-�����@:[�X�	����!�`�(i3,�˳�*C�����p���W�,�_sa��o���H�RtV�^����&��r��졾�g��]~ڣ]�,�F��P��}Dq�f����M$��2�w����� �.J�>��2�N�3����ۺ�u��ݚ�Н���w�w:�!�`�(i3��Aڬ&W�����=��w)��
=b~*��s�������P�íN=]b~*��s�������P�ڎC�?�M?��y�!�`�(i3����&��r��졾�g��]~ڣ]�<4�sg�!�`�(i3���M$��2�w����� �.J�>�u"����!�`�(i3�߆�p�h�	T����[�:
1���Ư����z��>!XM�#����+1�;�.��1�>!XM�#�=5.B��������xQ�1tSjv�!�`�(i3�o�t����w�`L�&�����~�G�kk�!�`�(i3ђw�)�WA�qIp��K/�k�2�]�u��y!�`�(i3��w�w:�!�`�(i3����&��r��졾�g��]~ڣ]���}��ݚ�Н��q�9�ͭ�Ƀ�?PA�g�+C��sJ�A7���ݚ�Н�fĉ>99��A0ok��
�:qEp�;�P�t�5!�`�(i3�k��M�h�
�G���69<Pk!�`�(i3&����aq���)P<�ܓ�Y!�`�(i3���4)c�ݘ<�̆x*��c�d����l��T���ӄ`^�Ad0t�;!��Q�����&G!�`�(i3�o�t����w�`L�&�����~�G�kk�!�`�(i3C�4M/�Sн3y��(|v��t����~=�L�~,�H�͛�!�`�(i3��\7�f�J0i�,�L z�P��*���k� �ԬQ����5��t�1tSjv�!�`�(i3@��( ���M/*�3�c�u��nu p��@���!�`�(i3i�:`�+PN#~8"�Z��q�����8���&�Ra])n#~x]V�{���>E-�N�Ӗ������%a t���~=�L���Z<��A!>!XM�#����+1�;�.��1��B� �b��!�`�(i3�o�t����w�`L�&�����~�G�kk�!�`�(i3C�4M/�Sн3y�ܣ{�j+���X8e��e
�:qEp'{w#/ B!�`�(i3]���\�x8�Q:��?��I�^$D�����v�)y�Eh�ѮYț��N�����*���k� �ԬQ����5��t�*���k� ֯���,mk��L�������&G!�`�(i3�7����������EN.�r6���`�v�l���"!�`�(i3ђw�)�WA�qIp��K/�k�2�n�)�� �g!�`�(i3�̢k���������PLm�<o���(4G��>� ��A�Y�
���3ʩ�V$=�b�������P�íN=]b~*��s�������P�꠼*d�m�'����u��r��!�`�(i3h5���=�t���_j������M���~�K���@�!�`�(i3T�=qއ*|X6و�cµ���(A�,"T�z�D�R!�`�(i36�B��~ ��A�Y�
���3ʩ�V$=�b�������P�íN=]I�^$D���������P�꠼*d�m<���H�
nЯ�O�!�`�(i38�_?��N�Cٺ����J����
%�6W����!�qg�L�[\�"��-����!�`�(i3�D�������{
B��e�g��%s����K!�`�(i3ђw�)�WA�qIp��K/�k�2�n�)�� �g!�`�(i3�̢k�����Tյ���#���n�W�G��!*���k� ֯���,�ۿ���L��0p�F!���~=�L�.ama�`m�>!XM�#�[��l�,t���H[W?a%��w�ݚ�Н���+�t2��Lq��QF[�Z9�+	�]
���7��*"(�6�F�}қ~�!�`�(i3T�=qއ*|X6و�cµ���(A�,"T�z�D�R!�`�(i36�B��~ ��A�Y�
���3ʩ�V$=�b�������PLm�<o�̱�	P �a��e�D.7�q���f�e���v[v%������=��w)��
=I/��\]� h�ҩ�!�`�(i3@��( ���M/*�3�c�u��nu p��@���!�`�(i3C�4M/�Sн3y�ܣ{�j+�f����It�!�`�(i3��jVѭ@!�`�(i3�D�������{
B��e�g��g!�%=F�=!�`�(i3���M$��2�w����� �.J�>��l8R��!�`�(i3HN��R��bP�63Z�t���%>�rGO�D mWN�ݓ�W����(�l9n�&U�)j�S<�6�Q=��\���S)M2B�FxU�?D�8�����vo� ��M�#�q9+t�}VA�ڦ�c4��Aڬ&W럼�~=�L�����3���'����u��r��!�`�(i3�<@���ل=����h����3��[<�m��I�!�`�(i3�J�g�*����3��?�4V�I~$�}>����=@'ѥ��Ra])n#]���\�x8��'��b~*��s�������P�íN=]a��o���H�RtV�^����&��r��졾�g��]~ڣ]�,�F��P��}Dq�f����M$��2�w����� �.J�>1�Ѯ�a�!�`�(i3�k��^�1�є��g��h�ѮYț��N�����*���k� ]�Լ�c�#o�]�ʄ�
%�6W���N�Cٺ�������u��r��!�`�(i3�<@���ل=����h����3��[<�m��I�!�`�(i3�J�g�*����3���˙�6Ï㜯}Dq�f��	��x��ݚ�Н��H�����K��I/b�W�
�rP&��dGL�F�z�>�/�O8���6���no;�M������P�íN=]b~*��s�������P�꠼*d�m�'����$����թduP���2�:
1����e���N�ScM?��y�!�`�(i3����&��r��졾�g��]~ڣ]�<4�sg�!�`�(i3���M$��2�w����� �.J�>�u"����!�`�(i3�߆�p�h�T���ӄb�3�旅Va�ir���J�sy�V��RkB�����X
%�6W���N�Cٺ��#o�]�ʄ�
%�6W����!�qgy�`��vN1tSjv�!�`�(i3�o�t����w�`L���$5� ����:N!�`�(i3C�4M/�Sн3y�ܣ{�j+�j)����r^!�`�(i3��i��:q����J�sy�V��RkB�����X
%�6W���N�Cٺ��}2��L��v��&�B
%�6W����!�qg�L�[\�"��X� 2!�`�(i3E~X�J��
�M���1F#�֞qduP���2�:
1���Ư����z���B� �b��!�`�(i3�7����������EN.�r6���`�k_�a)!�`�(i3���M$��2�w����� �.J�>�u"����!�`�(i3�߆�p�h�M���yt7�o�*H��& ��0>!XM�#�[��l�,t���H[W?����z����K��I/b�W�
���:�������7�|���޵.��gWaU �IH�RtV�^!�`�(i3�<@���ل=����h�s��m�Eq��}�[��!�`�(i3!�`�(i3!�`�(i3�qm>C`�ݚ�Н��q�9�ͭ�Ƀ�?PA�g�+C��sJ�A7���ݚ�Н��Ra])n#~x]V�{���>E-�N�&Cd�c��aj�\�T�g�����c��*���k� �ԬQ����5��t�*���k� ֯���,mk��L��x{^4��*m!�`�(i3����&��r��졾�g��]~ڣ]�,�F��P��}Dq�f�!�`�(i3�J�g�*����3����B����i��}Dq�f�՝� s�#���k$ !�`�(i3@��( ���M/*�3�c�u��nu p��@���!�`�(i3C�4M/�Sн3y�ܣ{�j+���X8e��e!�`�(i3���F��O��ݚ�Н�$f��_Ub����pT�G�&ց�*��JY�����ݚ�Н�
̛�]���n���G΂zG�_h�!�`�(i3@v��e��~$�}>���w�q���_�mS8<�n�ݚ�Н��7����������EN.�r6���`������ݚ�Н�ђw�)�WA�qIp��K/�k�2�������P9�C�s�4!�`�(i3�����!�`�(i3���g!h!���7�|���޵.�ۃVa�ir�K��I/��0�|섃Va�ir�K��I/,ܓh�,������&G!�`�(i3�7����������EN.�r6���`�v�l���"!�`�(i3ђw�)�WA�qIp��K/�k�2�n�)�� �g!�`�(i3�̢k���8�_?��N�Cٺ��#o�]�ʄ�
%�6W��M*QfY�"ZgWaU �IH�RtV�^!�`�(i3�<@���ل=����h����3��[<�m��I�!�`�(i3T�=qއ*|X6و�cµ���(A�,"��C&��!�`�(i31���~!�`�(i3�o�t����w�`L�&�����~�T7u��2�!�`�(i3:)!�1%�@�	^���yCw�Hm��!�>!��!�`�(i3��Ě�����}Dq�f�HN��R��bP�63Z�tG�&ց�*�3QAZ
0��3��Y$�M`�K)��v�:�-22�v%��v��!�`�(i3,�˳�*C�����p���W�,�_sa��o���H�RtV�^����&��r��졾�g��]~ڣ]�,�F��P��}Dq�f����M$��2�w����� �.J�>��2�N�3����ۺ�u��ݚ�Н���w�w:�!�`�(i3��Aڬ&W�����=��w)��
=b~*��s�������P�íN=]b~*��s�������P�ڎC�?�M?��y�!�`�(i3����&��r��졾�g��]~ڣ]�<4�sg�!�`�(i3���M$��2�w����� �.J�>�u"����!�`�(i3�߆�p�h�	T����[�:
1���Ư����z��>!XM�#����+1�;�.��1�>!XM�#�=5.B��������xQ�1tSjv�!�`�(i3�o�t����w�`L�&�����~�G�kk�!�`�(i3ђw�)�WA�qIp��K/�k�2�]�u��y!�`�(i3��w�w:�!�`�(i3����&��r��졾�g��]~ڣ]���}��ݚ�Н��q�9�ͭ�Ƀ�?PA�g�+C��sJ�A7���ݚ�Н�fĉ>99��A0ok��
�:qEp�;�P�t�5��6��V(pyL0D?yz��������[j?�{�X�[�g�DPp���ܐ�}��B7�Q�+ż٧����|�X$4Ƕ�W�S竚��ٓ]M\I��A$�P��O�@י����z��q�`���φ��<�6�af��pD���|#HK�����qD��=a�^7�1tSjv������ya�E�Rq���my$�N��o�/���;!�`�(i3+��/�6�.ZclZ�V���{S'���߆�p�hؽ!�M��9�a>*<UB3 �~k�%����ZAL�:.�
9� ���(ٗ.;���JTv���H�����pAy����~G����������&G!�`�(i3�'�c��dN�<@Iv��nt=:��:5A��p��w�w:�!�`�(i3/n��G�N_������ \L�1tSjv�<�6�Q=���3%�|�CH8W	ܷ�4D�P�S �9���1tSjv�#�աl��`�un�&	ܷ�4D�P��Z�I�u��r���&d,4���H��̣��@#('�cH_����d�b��w�w:�!�`�(i3��$F@S�� 63�镋�%>%��
�:qEp�;�P�t�5����l��Ϭ�g�(���WxdZ#'��� h�ҩ�!�`�(i3��Bf���.��!wx�F���m¡
�:qEp'{w#/ B!�`�(i3��NƥN��nF���<�W�.�P�	��
�Q�}!�`�(i3�5ߧE4��!�`�(i3`���*1
�:qEp�;�P�t�5
�:qEp�;�P�t�5fĉ>99��A0ok�׹�F�}�WP'����~͏/w1z��ӊo�*H��&Vi��pb��H��̣���ڻC�i�;��|B
5�v�O?�d���&����r�6/6$�S�1���L���|��Ծ��i3a��o��_�Rv�䩲$����E)e|A��`���φ��<�6��7�癆cgR������������ h�ҩΪ�\���S)k	䶙%T7u��2��k��^�1Aj��t�35L��$
8��2�ֈe1tSjv��o�t���Y��@��( ���M/*�3��E�i�m}6O�D mWN��ܐ�}��B7�Q� )ZX�B,��ف�ׂ��3�Z�#a���_Vh`�����!6�o8:4�I���c�90Mj�dL�{y����i�q,?5q}�P�|��U���e��d9=���u��r����3�Z�#atw�t����\��/.f1]�?����Ro�G/]%�z�-uͺ�s�η3G��Hb� h�ҩ�U�07�:��=����h�����$~@8c���L�Aɠ�T�nGHN��R���ء�I��߸��S�Ȍ^��,P�H����_Vh`����2g@��?u���\W��	]�	�U��)���Y;e�iK-pm!9�>��n4s1�U��B��-��^�uJ#��r$ɓǉ�.y�U=������&Gђw�)�WA�qIp��K����^7�j)����r^��$���͜P_�_S:g�RMm�o��'����u��r��T�=qއ*|�O=�W��K�VSƅ��	^���y����W���Ě���aT��3G4������4q0�I�ݡ��1���t}�F��<�3y�� e
)�*U�a�(���Ņ�F'φ��<�6�@a� ����C�'�ąd�G}%����3f�;�C�f��wFlE� ��'ž1�|��P�:k& 2�]�<Ęy��j��k$|�N
�`����;q��b+}y[^	QW�Q!r֯���,��e_cƍ2���l�J���hB;����� +��$�\%e��}Dq�f��K��I/��=����%��v�ڮ_��>νr�T�g�����Mt�꾸b+}y[�k��^�1��dc�@c�����h2�]�<Ęy��j��k$|�N
�`����;q�"��ӌ�r^	QW�Q!r֯���,og�Ѩb�����=�#����=ᜯ}Dq�f�g�G��0B����\�����$~@=7�7K�PO`�� \)������P�]Z����?�4V�I��1z�a���������~=�L��i
�i�w��2�N�3�`tuL���$f��_Ub���uQL+��φ��<�6�8���SY�N��&Y��V�@pن���v?�����觲��h�j;�U��)���Y;e�iK!���d.���+�^n=\f�5>�1x#0<-�1�}��u@:������r$ɓǃl[�Ƶ�1tSjv�s� ��<C?�����觌	�����e��0�U+�qbp@��߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#�hҜ�����!3�o�O��-�����_��>νr��U�,��/3�|* �����2�N�3�
R��?U���%>�rGO�D mWN��Ě���aT��3G�IX0F�M����S���G�M��#����'a��[��l�,'���R�+���7�|7�O�e�^��\���S)��)�
F�p�YD<=�������kOC����x�d��::T�����ևA��݁z^'���>;#9���Όe������P����A@�-��T��E�����y�"'�w���g�Dp��H�1!�J�G�~w���q��߲�1V�L�H�^A02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-���f�ӄw�c_B;����;��b�^"BL�|��{+&h��z#�|s�c��D
�=I���!�)¾�O�aIE���R����+��{"X��/��m
>c�.[K��m�n�Щ�[���(/��""�i����E�&�F�i�J���VKp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h��v�{�m�D���JG=yg�#w�6����#�W�G��!?�d���&��������?�d���&�τq"�;Ȋ��f�X�w�&�Ԋ&b��@�A�KRM�,!hޖ�A$�P������5d��n4s1�U��B��-3��܌o��%��q�����"sS<�0�zG����ZAL�:�@��v{�G��R:k�ڛ���Re�
ƍ2���l�M���r8��]�p� ��߆�p�h��d��JXl'�T��~��Uг�|<���vo��VF�˷��E��Pק�VF�˷���}Dq�f��G�-!�5/�V�q2_�mS8<�n)�{6�U��-��)'@�	}��Ԣ�"u�����`�����>}�U��4~!�`�(i3M���r8�Q�lՖ�?-O딈pᜯ}Dq�f��	��x��ݚ�Н�����������**,n����"�$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vx��e/1��!�?�����"ZD"m{�&�E�3tM��楱�o��_�Rv�䩲$���o�,�T�iI9�o«IX0F�M�����y�8D�r^�Hd\���F�`yx�>�+X�[�G���K�k��M�^���+| �Z�_v(��ƍ2���l�E����[�k�n�=���b+}y[�̢k���F�KD�Vr[/}>5��0jJ�_/�+�����l���n*�sL��.1x��w����֯���,-}���A�a��o���H�RtV�^E����[����>^17Ӿ�b+}y[��+�t2�4\%��t����{���}Dq�f�-��)'�	�;���x��N���!�`�(i3eX�LG�5:W�^�|�����NM������%>�rGO�D mWN����l��A�k�C�
�u� |�[��CC'ێ����� h�ҩ�`��v
K<߲�1V�L'�^�����ݚ�Н���Ě�����}Dq�f����F��O���\_qFgyO�D mWN�׹�)��, q�&�E�3�P�k�P}Z��E��3?�d���&���v�{�m�
�9��������F�U�S��5�����h^���门:<#�'	�?��[��ҽ���~���\�X@`u:j1�e�Ǧ���P�7� s�7F�S=B��{z�n�����s���K�A�'$�mo�6LD9�����w�R���y>��yС��P�Rn4��8L��!�`�(i3!�`�(i3!�`�(i3"WK�o9z��_�^�]_�ϋ�G)?�����s���K�A�'V�T_��p���q�sY4\%��t1~��;h�������(ݿ�O|���B��C8�4K��7� 05
������oA&��>�~q�z��µ�퇇М1J�a$�Y �����s���K�A�';�¬pX��g��U-�e�j
��z�Ƅ$�O���z�j�S�Ƀ�?PA �+�v�<�fm�oH�	^���y�,��z���:���05ǒ� 5T���Z'�����S�uG껺<�]iO��Oӕ g�|�a.�Ϡ|&����x��B�KS���H�	�k�~N꛺7&���LUFƗ\��Dz���T��/:[%=ѵ5��#��u��I'U� +iF�"�9Ϭ���/�MYN^�?��΃�����(��H~3%jA�L�� 5T��vb8��HM�"�5l����k"eK�$ϙRl�bș�� ԋ3�0zYc�[��F��S�J�w��|��$�5����Ou�X#*ݔ�	������3�Z�#aH����U��)��S��PL��=7�7K�PU���;}�F�e{iʖ.���0�v��n�ƫ�}<�g�G��0��أ��B�/N���F�W �{y����i�q,?5q�kpR,�y6�T�@�\���0�Uui����0�/N���7Ԝ7(u��ݓ�W���q�Eh�^(����K˖�sM`�K)��v�R�<<�U����$~@F�e{iʖ.%_����T�KKnf�܋�n焞	�Ȗ@@��H����g�G��0��'���C&b~*��s�/$�ߺ��]��pZ�ì1F#�֞qg��J�s��{��b�b�*������� h�ҩΖ7������8R ���M/*�3�2�:�#LA������� $�]n�ݚ�Н�T+���fS�n�(�a�:91�7ՃVa�ir[��l�,1B��CSk#o�]�ʄ�ݟ�e/�dI{�8k��.ͥ�H�RtV�^�D�����0	�+G�c��=����h���6����'�I�َG���:^E��߆�p�hب�������kO�d��-��!g��J�s��F�e{iʖ.��4�JCk�!*��*8����Uy�`��vN1tSjv���+�t2�;�������w�`L���JeJ��5�W��@�A٪�o�_&�
�:qEp'{w#/ B����&�� ��\�&ɖ��_j��� �5�������m�Qfĉ>99��A0ok��(*�O�q�Y�G���֗*����ْA5��9�O��F���R:k�ڛ4a��|�&��}Dq�f�}I�6������U5C��r��&�����&G!�`�(i3U�07�:�tMɶ���74/����G🕾{!�`�(i31���~��+�t2�;�������w�`L���JeJ��5�W��@�Aw��1���.�\��$�$f��_Ub�F�S�1 �����$�W��@�A�a����I��ݚ�Н��K�,ǆ�`�܋�n焞}��NY��}��-����!�`�(i3�,�B���{
Bg2�I�7�js�і��D!�`�(i3#l'U:�g[-�¾L���I����~u���NM����Ra])n#���r�����D�����0	�+G�c��=����h���6����'�I�َG���:^E�����vo��VF�˷�!�`�(i3��$�\%e��}Dq�f���Ě�����}Dq�f�� ��F�	kwJ�Rmv&&�6,d0AL(�z��?�t�ϗφ��<�6�U�07�:�>��1]��a� ˭M�ʕ�I���܍,6��zU��'�¹ӱ�_r�e~5�O�%E#P��èV��d.q��9�w��H[�Wi�(5���2������<�b�5L�T!t���m l�o66����~�����!�sY�N��}�kmPک>=�[b.N�ؾ?u�^���_sM�u�2�4�*�s)l໶�, e8�~����U���a~�'�� 7��
�+�0ݿ����j&�>=�[b.���9M�o^���_sM�u�2�4�*�e4���F[�l�e�'�$Zյ[+8�a�)��Ƃ~6T���Q�x1�~g_�,\ަ�It��+g[�Zt%��m&<>��%��JU�a�(�n����62�tϛA^��'T���+M�Mb�:u�w�vG�q�:�&����#|�1�0j��*������Э~���V��2
L.�X;p`��vbëdP�4e���>�f�?ǉ�=�1_�
774\51�]2�t��MJT��
!�7�R�"�*}#2\z��``�ǆ�!�`�(i3�&8�,�aG�	�AS3f���])ܟ�Ma`_��r����N�i-9�}�~���lscX{�X!,!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�;�
Ơ�*�6�M)w6(��.�����gRI/!�`�(i3�Y�M����4Wt#��5Z���r����ؾ<k�[��x�ܽ���X;p`�T���'/�>#2\z���&�3Z�K�!�`�(i3�&8�,��y��ЉT�9e��/�7�(��.��?�!�`�(i3t$Q���V�T_��p�V;�������gL�4�2s��2 !�`�(i3��5@~JuM�D���!�`�(i3W�4�:*n~�<�&��Xh�hk��a��OY�P�CQ��Bރ;�{��C�{����K�7��(�mWƒ�a�}�$Ϩ�;?���*/�|�-���w�E�V{�!�`�(i3�;���5!�`�(i3!�`�(i3�<��N�L!�`�(i3\��p��i�6������uSKA��g]�RN�]�5'p����nZ���t��˳3[�u8�|�秽m-��#l'U:�g[q�vG+|�<竷b��"&�_~�:N�t�%�Z?��<�ry^�C$mQ���&8�,�(]ͅ�y�����&FM���hy��jX�p!C+H��bf�?ǉ�=
���&~^)-�����4)cq�vG+|�<?V��j�cc����L�{czZ�����f��8�H�ݚ�Н�*��^�"~H��
�[�<�`A��_i¼\K��X�o|3xD�̯ƭU8�$��`���	(��7��F�dHP����|�J���-M+����"X��[O+oF��}�;��������/s9S��I�����Y>�څIׇӭ��*��^�"~H�*�qAW�j���H�D�6U��OM�ݚ�Н��AO �X;p`�B��C8�4gG��M�ѱ�ԕaOf���x�f7﹏S��I���f�E�7��RN�]�5'��t1?������V?����(sW���4���M�{�|L���\:g��V����f ���t����G��F�/L!�J���B4�@	�u�a�ݚ�Н�!�`�(i3!�`�(i3!�`�(i3��kw�G�I��)���W�w��fD�:J.]p��5�!�`�(i3!�`�(i3!�`�(i3m�ڨ�hծ��d.q���x�_#>����(gR� �ұ+s�Di�R{LdR�?�9�e�D�a~�'�� 9LX��O2��,���C���:4.Wr2��B���z����^�~����U 1�|�I� KY�!�sY�N������?Z~a���@=�y�z�5J1d��+r2��B���z�����\�Wd�U 1�|u)W~ۚ��5�O�%E#P!�`�(i3!�`�(i3!�`�(i3� �i���(&�L����K1�dѤЭ���PM�^-q�x�l��1:�N�*�xSƏw0�����*0e�El����ؑ���6�M���ʄ�F{/����MB�8"FeIN"�-���0�i.�9Ɏ�#���?���,�v�q0�~��̚Y�M����4Wt#꫕��!N �ݚ�Н��L�K��%<7�`+Al��R��������,NL ���X:��+�<6��$)K!�`�(i3-��iW��
�!V�ځ����M���7>���JU����^b4b�;��Z��i�ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3w4�4a0E5' �c�X�0���X�q!�`�(i3XO����0J�y��*?(���6%�a(��.��/��lӹ��zigzA=v)���K�7��(�mWƒX:��+�S�9;/���!�`�(i3-���j_�ܘP{ǣ©��,3�/�r^w��'�k�f!�`�(i3 �R!�xY���ݪ�7��?�� @:d;=�hKV/�g#2\z��}�� �с�'(�U�c�&8�,��
�Q!}-[��u����g�&�0mB7Ԅ��7V���s�������"�9(��M����v�v��8<e(�y�|����x��~iM5/�S3 <�X;p`�T���'/�>X�o|3ԁ���T!�`�(i3�&8�,����0u�C!�`�(i3�g� a){��Rk��?��q�M�4�a8&N C^�e S]#�e����kn4@Q�/�!�`�(i3 ��$�,����/ӳx��R:k�ڛgf�mk�X�ϣޓ��&8�,������	�;�ݚ�Н�;7hZWT��X;p`��m�Euk�jB,�<fI,�ttT��Q�#<4^����*[UxG!�`�(i3~n���,a��/ӳx���{L,8gf�mk�Y�ay}M��&8�,�6.���͈�S;��ܺL���'T���+��PJU���ӊ�8�5�Щ��O�*���]�ܯ�Կ���p�]K&sӇczZ����/�e��<��(���B��������R�!��+�g��U-�ew�K�H/��l\�6�'����7Z��$�~c/z��q���P�;�/O�M�Mb�:u�!����3���3E M0�~�O�������؟O�!�`�(i38�$��`��x�i8B2�GW��*���i�\!�`�(i3�$�~c/v��&EA)<�!�d�<�@O��YY��_�,)ȍHK�ZHOh#��ڥ����Ⱦ����G9L�M�7��<�vW4��`�}d�ȢiLO�����=l���d��F*�L��!�`�(i3!�`�(i3!�`�(i3���D4FFG .٤��	w�R���y�A[�;���eF|YTF^�T�r����!�`�(i3!�`�(i3!�`�(i3(�JZ�Vk�;��|BI�]�,t�x���}���_�T�:`�\.�IbR�K���s��$�Z;��|B��� OD=����Vʆ7���өqa�*���zL͊�q���c<53?���?#��4�Ց�ʁ�X�W��vbëdP�"��:b`��/�XD��(�[6L�}�}��<�ԗ&x�#r�����èVp��E|��t���7�I�?g�f%��h,��;�0��'>_$MTy��9����S���� "5�]ޥ0D���3A�)Oq�i�-}�[�����U4 :��	��aJ �!,P�H@��&-���xԞ�����i��E����p��x.�Knq,���9^-���2��̪U��֜��3�&8�,�e*���	&���`"�G����?�s!�6]��E[WͶ
�`��~mi�ݚ�Н�EfVNN�0|]<w:��X;p`�U9����u���q����k��,��C:���2��}��=�lx+~�S��I���i9>���Ef�?ǉ�=�� ߌ��-��Vi� �Z�xOQ��B�'��a���p��b����z1]�xv�:��p=�n�Ԓ��K�u�c�$�~c/���F�ƻ!�`�(i3~n���,a��/ӳx���{L,8gf�mk���b~y� ��&8�,��Om�"���^���F{/�����,([�y���㋞9�nX�8j
Jt��)���l\�6�'����7Z��$�~c/~�O�������+�t2��ӱ}�tMTl�����)��.��f�?ǉ�=�M�g����-����b=��y��j��k�lԇ�-{�4�0 L?�p���@Z�6[��u�V�<�nbBIճ��)��]m�(�h@)í�_�ߍj�������� 63��p�@OM.IrP"G�wk��jr�!�������,\������,Y�I��/^�=O{Ue��*�̞��>��vbëdP�D�R��	ܷ�4D�P���I`���jVѭ@!�`�(i3!�`�(i3!�`�(i3��7I���
�)W8��V��	��y�㘞������8I��2�HF�M]y��Z�/�N���N
k��L����4��>���O6�o8:4�I���c�90Mj�dL�{y����i�q,?5q��N��)�Q��l�'ž1�|��P�:k& ��-�����D������"r�V�)P<�ܓ�Y�̢k���F�KD�Vr[/}>5��0�B� �b�Ж7�����5*A�u�������$~@l����*��"���l<o�;)�y���ƚ_��}�	76�&�� Ӗ�t$�)�vx.F<!W���zՇK����3Ah	)ޟ-�b�+�