��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�~09h�i�Nq�{5��]�0�lK'���Xw����Q4?���ʢ\��|�����o�3t��v'gn�]o��in�m��+D(m.�B����s����Ct�z&��ÃlO ܅doGa�젿��ʐx�?WA{I�Z�T�����N\� n��A�T�g�v�;�K7���'n�^0o�)�?�^�?�XW������w
��ڎ:�ڛ)
�}��ɣ�YV�PD�E${��4`�˨�;O8�d�
~�n�}Y�:]�@�<g��ũ,+$\�M��lJY�Pt���`��8��f�`��[��Yt��'�d"[~6����aD6&>��Y��q��f�}��`<Y��sp�����5	���]���c�A�L'�������W��_�ړ8���/��4��}�<�N컽kg����|g�Y�'���Xw�j�7����'�e���"j���b7|#9���Y��
�iC�E����F��j��\w��0]%��C���+�
�c�~��j��\w��0]��0�&�ͭ�E����F��j��\w��0]{k�h�+m��q'��7G#+�Ǘ0z�cUL
 '&1���D���J��8���/��-�
�]o��in�m��+D(m.�B���B+F�bh������R(��z�jv .
L����1�:�Ω�`��G��l&K[�
C�m��P��I��'�Po�Q�>�������IÙ=�HAmY�f��Ea�8Ss�LPo��p�(�oE��(��f��Q�m��'A>􏄃'�wZp�m~|��SpX�@>׼�\�v����ř�L�g?_��<'P��!jcCA�T�g�v����fQf��p�m~|����F}x�JHn��z�y���݈eG��{Ǧ%W& s���r7�����^���I���P4ǲ ���h9�5�܈zc��%��XP����c8?-+eN�Ȅ�4b�rS�b�8Z���'�e�����"�?;(��j67�Qs{ɯk�>p�m~|��7�q^�1�0M�/�s���'n�^0oy��\���W#�i'�6:	�<�&IMdK�Ch��T:���V�S�ff�݃зq8�Ј'���Xw�j�7��Po�Q�>°������R�wX��}�
�?�`<Y��sp4�r�@E�n`5�fK��0z�cULn�4Z_U���l�����"X��[��Q[R�7����n9읖w�x�z�f.�Э]�d�٣��c�A�L'�"��/f~�ƃ
ᾆ�x�T�\ ��i3�|)sՀ�T:���V����̵?oзq8�Ј'���Xw�j�7����;1�˚���ӯIJ ��`y����@����gG�������+N�f�+��Q]� _�rs�i�76b�*Ғ�ߨ�,R��g��U-�e,%�0g���l������*b��93��bj����Z鎬�������(������oD2��Я�R�wX��}�
�?�<��0n|�!h�b���t5a�l��0z�cULn�4Z_U���l����g��U-�e�ˍ[L/}�t%>^�ߒ.�qO���WS���
���A����|�������-�YM*b��93��bj����kѶ���� >�������.�Ӂv��9Kd��"�����ڗ�\���V2���<�؊�"�Dz�Q��y{y����x��F�U| c�]h��)�MUK�>K���T7���?kg�w�4�ksĶߨ�,R���"X��[��Q[R�7!-B=�6f1_!��Xm�[�̷��3h��;1�˚z����'6���;8=�g��U-�ePo�Q�>��Q������w�x�z��!�L����� �#7ۏs|�L;Л��|#9���2jɸ'�L\�z�´��2jɸ����oD�O���j����k��$a(􆿳���GFwk�ߝ�s�P|~-�6ώ�<�"��v�aφ��<�6�@a� ���N��ȥ�n4s1�U��B��-V���$��bŋ~���%.��D����A(�c���_G��Hb�8�u?��I!�`�(i3�d���a؅q$��.��m�f.���G�?v��� �+��R��?V��j�c�ШT�7VE�g�������(ӈ���m�r����*qA����6\�4�@�� �-jېI�q������ л��E�BS�+��U�,�P!6���r����L�J)���� \L�1tSjv��H����!�P{� ܄��w�J�WJ:�f�a��o���H�RtV�^q�\E��0,"�-�˺o_B�E�JX�Ή������$�����&�%������k��$a(􆿳����^��Ra])n#���r����q�\E��0,"�-�˺o_B�E�JQm��	����$�����&�%������k��$a(􆿳����^��fĉ>99��A0ok��$f��_Ub��7��G_���;�P�t�5�׹�V���$��bŋ~���%.dX��҄=Z��	�`DÜk�K��h̷_��yC��S8�\�w�4�*)�2�"ղ]�6��2�~�P��qa���=7�;-�]����2jɸ]�غ��>���f�RE3-	�����3�#��rY�{'%s��$��S���b�Bϱ�!-B=�6f<Q�vn��l����I�/=k��T�'Y��P�RG�;!�`�(i3!�`�(i3!�`�(i3!�`�(i3h큈��]v1�_ُ%�W�%�KY��{&���'6���;8=� ��g�SE���̵?oJ�
�����WYHp(�e�	�<���!���c�A�L'�ɻ�L�1p/-��ս�9�j�����oD�d5z�R��5 �8��B�;j!%�)��=���!�`�(i3!�`�(i3!�`�(i3!�`�(i3P"G�wk�Z�d-�~Ee�1���1�����b��[� p�!#��Rh���K�6���!�`�(i3!�`�(i3!�`�(i3!�`�(i3�(]:�z.��Q���_2��VU(��z�j�6f�L��.