��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�"� r����`,��I�|��]��;�Iώx�t���E�L#uc��WŬ�+�-ޗ(huUPc�k�u�}�R�6�_(!��?��Xm��+�����l&K[�
CN<��;��� B]�pE���	x]̃Dj#^Da����M�r���
�'�ө-$J�z����)�,�˛D��w���旴4�����:��@���b���$[G��m$�;�`��v��p�㈍x���t�켻�S���c,31�-elwB(�93;2���Zߧl4���0�?�1~�x�c�>j����d��S�W�>��Q�d����t�mR��:�����-��3���7�Jk�b#Ӡe��?�F��&��q�©�����[��&�u�"��U���T�����\�4�slom��Q�N�5�%W0�ր� !�zA>(!�o@���q�&2�Z���8fw��[#M����4L"���ې����~I���&���M�|(Q\��(��~��I(K�b	+��~ķDh�D.�1o�����.��:o(~'�@
��,:�Y�ͩ�,�~�B[��Th_&^�� �T�9�Y��6��X ����W)d�H��K��Ap���`"�E+�-_���^*s&QL���BPJ�%�9
Xߞ���������b֡�0��RL�a)'r�Ӟh� ���G�/9{�d���D
���PJ�\�����A�p
˽0?�.���*��� 9ٞM���]��8����t2�}G	p��#}�{�Sc-@G	>��RL�a)��F>x���,�%���pY�� e��x-����l�;H������K#Q�����1�%1�����:�
�~�K�K^Gc7/��#j��;�i1�璠�J�*��f�I��r�O��C��0���۞�^��u�?�L���zZ�Y���;H������K#Q�����1�%1���
�׺R}	C���`'�t?��<6���'�t��,l����k�8���҆�|n��T�{ ��ʥB�2��;��u���^G`J�Й�m��/K5r��!����%�[[e���|���>�
� �AH�*��.�T�{ ��ʥf�nm��mHG���i�P�Gy#����*��jr�4��X	�ƒ��c�w�A��P
T�]���X����PIIN��d�=o����"���	x]̕%�h�Gqc�J�M=
�ٽi"���g�aa�y���bAg�
d�m��+����o5��6V�|��f$ui�V�3ޕ�L��՛�;��4�W�]�a5��6V�|X40��7��XݓAA����~�9�؇�M.9$o��݉�X��R��
�A�`5��\�4�si�W���Y��݅ 00b�������x�o@���q�&ϖe��!���q�L���Q����m�!=�y����h�}���Hے�8Y�&�\�M�C�вC��J�/�_?�hbHp|����#�n�%@ܣ���m2�5�A�E'���M�Պ�s{�tA�~�u��,6o�-��ΐ�?��A�}n���t�o "�xCo9�Z�.�"�K����	x]�G�Lm=�b�7��Mv�9]Sh��3a��$����aa�y����>�u��8#t����nr�O��C��0����"g�����I��s���1�#���Z��\�����Og����n�&\�ƺ���m�!=�y����h�})6D�T��8Y�&�\���
���;Ppo�6�$�PT8��Ì{����V3��p��b��g�|h�03�
� �AH�*��.㤚{y�ڵ�o!f��L_!�pN��i�P�GyϪ+2�Ľ��3rn{����V���	x]�<���e��8�t�~��,�O�W��s�!5�S��H���)��������ҥ{E�?HF��eUٻo���mi��*	�ť�.^�i��' 1wH�x�xs��3�<A��z����
a�������~�+��,/,����W >g1�]l�&Y��F}갨y�����# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��`y��f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�}�Z���ik2)�
}wʭU&H�1��8�h7H�u�ÍeRuw�C?3d,f$�7Q0�"<�F�ٴB�I�SbW9�v�H�F?t�)�Y¹w�.� -��E�I�?g�f�Jm*)�m��+���%	v3l&K[�
CQk�� h��ߖ�g��o�4��?����DNZ�j׫���?_W�\I��ఽ��`g�5��!08��r����N{a�9O����T-Q3�Y	���,�V`t�iZ]XF�������̅�ԜF��v���N��!�`�(i3,ԯ���gn�yZ��͠4?:��X��yM��#s{��'�!�`�(i3jݭ�F����K������]V�H7'�R�^Ƒ��!�`�(i3�E����F�Z�>)��p40�zɈ��:��W��?5���{�z.�]�\�Y%T��BP��&��J�1�KB|1<\EfVNN�0|]<w:�!�`�(i3=]A��O�T=�4e=��-�ĕ|G�������{������T�κ��Cj���P��5B}�=Ll���ms6��	�؍��R��j�.(Wx*�ꢤ�OgB�Y���c��|g�Y�'���Xw�j�7��ct�:��RE��W��_�ړ8���/��4��}�<������K�]2�y�Z鎬�������(���`$�P.eE���lC��U�T�\ �͹g}|�H���p��b��e������]�!��	Ǹ�y85�B���0���^̽1��R��ӟ-�F`���G���`y����d�cCKA�lG�zv!π�����
L'���Xw�j�7����w�K�})9ͬ果��S�<Ԣ�7Z�:1�\mdЧ^{�j��$�'	����Øf� ly����)�{� �"c��Et��q���U��ͬ�	A�/ї:��|g�Y�'���Xwem�B0赓,([�y�|���(Z鎬����F�71�B��0���Y$�Yl���#�]�!����M[��ǢJ*�8�P:�����5	���]���>����C�h�'f RY%T��BPe.��xu	�>��l%i�-̇i�d�?��E����F��j��\w��0]%��C���M��cg�P��-��%M(0̈��N���N�?�_u�-����#u����T-Q3�Y��x5	+�ˬ>P�2-i_���F�� �yz��$6�.r-����G��9tf<[��H��֤�7ޚY㮭����t����g����=JHn��z��x�f7﹏!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3��p˪{��yM�B(p`D҉̖�7�j2��$q�$�È�P4ǲ �U�W
8�[q�<�J�G����\�v�!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�����籎�ʹ�q鋃+�y�^v�;���p�m~|��t���A�X
i��t��y��Fp����f���,(���B��ɓ�~Ҡ	��[�)�D#���ߔk�V\�5��|�~���ł�!r�97��EN�t�
�l���yM�B(p`D҉̖�7�j2�ف������̞��>���ԜF�����`���W�L�sQ������f�k� ��]�}�
�?��#}�{�@�m�W#�����O�BP"G�wk�١��	;q��^̽1��R��ӟ-�F`���G���`y����@����gG59#�X+�ez8�US�б �A	�xZ��j�
�iB{�Z�_��㶢�&-���x�F`���G���`y���h}Nw��諚��y�[�9=l7�kD�]�!��	Ǹ�y85�B���0���^̽1��R��ӟ-�D�s�A6�&-���x���h;C	�T�\ ��i3�|)sՀ*�şxˏ12v.^࣡NxZ��j�
�iB{�Z�_��?� Zh�RG�p�P�"i<,��1��yM�׶��	��:�g��U-�e,%�0g����Ed��>�^w�=�J�5q��T�ٮ|�,
���A�;�֋`N��7�j2��'Kb�|n���7���ө�O6�]Η^a(􆿳���2����.〧I���>G�g�����K�M�{�0z�cULd�g>57<�C�u)�6�3A�)Oq�fhz���I�Ūeߋ٣�o{�i7�v�ԯ��Q[R�7��s=q�SJ;_Q���Q�����&/�\[$Q��
�̞��>���I�Ūe�ǩ"�4s2��ԜF��g.�~R�(�%�8�ټ*w2�56d�x� �q��Αk�]I	V��@��/xZ��j�
�<�rם4�SR�wX��}�
�?�����E�El~pDa�G,�A@��}�Y�ןw�8���/�I����"�����,.��J�����E����FZ鎬������_�,��)׺������U�� ���E����FZ鎬������_�,�ݫ,��G!�`�(i3�E����FZ鎬������_�,�i"��n}n!�`�(i3�E����FZ鎬������_�,���o\<��m�HT�AY�E����FZ鎬������_�,��T:���V��c.��V�E����FZ鎬�������(���`$�P.eE���lC��U�T�\ ��i3�|)sՀ�T:���V��Kk
�&1�E����FZ鎬�������(���`$�P.eE���lC��U�T�\ ��i3�|)sՀ�T:���V��^7}�X5�E����FZ鎬�������(���`$�P.eE���lC��U�T�\ ��i3�|)sՀ�|[p2e�F;p�	���&Ũ�Z鎬�������(����F�dHZ�F�\Ȳ�r�r%)cA�z���a�R�wX�ո@����gG�!��V�B�b�Xϋ?@7s�9���o��S8�/ #O�)R�^Ƒ����"X��[��Q[R�7He�-�c��e��Y֡���t���ό���.�}�
�?�L�ԸK�F��	�c;�Q'���Xw��
IǬ�9PWC��ٯ����!�`�(i3��AU�D)y�Q\�@vs""��Fq/�bi��;��|B<&ǒ8�|s�g*n{��)V��B�1'���5�d�cCKA��0^˥�2��Gg�5rU�U��)���Y;e�iKI/B޾PԐ#��go`iI9�o«IX0F�M�����n��
/��y;�!�I=�+���r$ɓǃl[�Ƶ��I�q����!�`�(i3�d���a؅q$��.��m�f.���G�?v��� �+��R��X�o|3J;_Q���Qs��>H�,b�z'hۉ)S���o�Ra])n#���^a�nu4Bޗ��jw�	�����y��lD�7m�T��Ʈ+ˀa��z��2�,�s�Yls�<Ԍj��_�mS8<�n�ݚ�Н����^Kho�7�j�Γ��-����!�`�(i397*�SCj����I~E�g�������(ӈ���m�r����
�:qEp'{w#/ B!�`�(i3���ifz�d=+ӓ��#!�`�(i3*�˜	���x�Z��x�x{^4��*m!�`�(i3;�jmT�#-����p������h�'T��x.�Knqd��^��R��ӟ-�~�{ ���ݚ�Н�!�`�(i3�Lt���h%�㱰�!�M3����k�����-4�{>��!�`�(i3��Ě�����}Dq�f����%>�rGO�D mWN!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��jZ$��k�4��x�S~p�A�W/��WuV�ǵl�j6j�"Hs�����/I�|w��!�r
�ޮw�`g^i���E����FnA����hy�Q\�@vs""��Fq/�bi��;��|B<&ǒ8�|s�g*n{��)V��B�1���k�}���L�B��HJ;_Q���Q�X�G[��ht��R����A$�P������5d�`UNP�{y����i�q,?5q�c^����24����S������"sS<�0�zG����ZAL�:!�`�(i3�� л�4�>������9�@f���ʦ�/\<���tݻ�ݚ�Н��Lt���h���pb���e��0�U+�qbp@��;b�-�2�k+Q�h'�Ȝx�5W ��̫(�8�u?��IlG%��`��ǚ��ظ
��@�U#;�jmT�#��"����G��Hb� h�ҩ��H�������bO��M?��y�!�`�(i3p=�n��jP&}�mdN�<@Iv��nt=:��:5A��p�Ra])n#�V���p���y��lDQ�26�'��'r=I4�!�`�(i3&��f�_"	9צurT��âh�{~1JS�K{a%��w�ݚ�Н����y��lD�����
��.�)�p�!�`�(i3��ށ��yL��.1��\��~UD�Xy����I/��\]� h�ҩ�!�`�(i3���ER�.0R��崰�7���ө�)�F��3A�)Oq��r�۫�a q��j�J^!�`�(i3$��yx����WQK��<�7���ө�)�F��3A�)Oq��r�۫�a q��j�J^!�`�(i3$��yx�����:�z���7���ө�)�F��3A�)Oq��r�۫�a q��j�J^!�`�(i3��'T/��2������M��U��w6Q,���ʓ��m��Ed�c�B� �b��!�`�(i3X�o|3J;_Q���Q�=8Yø�Ӆ��g�Bp�>%���-ǫɒ�!�`�(i3fĉ>99��A0ok��!�`�(i3��i��:q�5/�V�q2����*�
Z�y��	����VPYu��r��!�`�(i397*�SCE7��"�=r,/��g�ŕ������!�`�(i3�	��x��ݚ�Н�����l��A·�a���ڌ�&-���x�'@�(��P�G�p�PB��r~�!�`�(i3!�`�(i3����P`��'5Tde�أ&-���x�'@�(��P�G�p�PB��r~�!�`�(i3!�`�(i3����P`���-��Y��&-���x�'@�(��P�G�p�PB��r~�!�`�(i3!�`�(i3�QX��?D#�k��5:�'��k�	6��J���뇏n|,�R1tSjv�!�`�(i3�Կ���p5��6V�|q��c�3�C: ߏ������'��p��!�`�(i3fĉ>99��A0ok��!�`�(i3���F��O��ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6��Lt���hm�(��k8�ڶu�7�w�R���y�Z��T�.�a=�J�*;;�`�D��ݪ�-oc���u�(� rRN�qD���o��_�Rv�䩲$���dS@Ɵ�o{y����i�q,?5q o�n�J-�X�G[�%��<� xjzӝ���I(͂�'�ɳ��!�`�(i3<�6�Q=��S<����K��!L��3w #�T�Z��&�2�����kv޶Gl�e���;���
`_�,\��ݮc7��h��w�K����+��dЧ^{�j��v�9��rI�F����ez8�US�б �A	�h��,���ANʂ��t�Ǌ,6KX�#���x.�Knq�n��I[�t��#�Β �r��!�`�(i3�^E4+у��b�Bϱ���ԜF���v!��c���w�K����+��dЧ^{�j$��XCp=8�b(��Xo=��-K��y��j��k�����5��"'��e�(ŧƇ��j)����r^t�R!ME�б �A	�!�`�(i3'�^����b�0"qo�0�ʂ�j�Ï��	�l�lM�3 zM#��m����F�P�7��S��h��d\��H����o�γ�ha��o���H�RtV�^�I�K�B(�W ���t�1tSjv��B�'��a���p��b���ez8�US������`�K7͍��|��W&":�ݚ�Н�f���8�6�e���;��U�� ���^E4+у��b�Bϱ��MQ�'����㶢�&-���xԲ�Z��*�!�`�(i3�5?�&P-ߑ����������;q�,\���q���7G�p�PhaWr��ڂC�u)�6�3A�)Oq�fhz���I�Ūeߋ٣�o{�i����zf��/��@���-��(�Ļ4��aA�'�I����~u!�>!��!�`�(i3��v� 8�e���b�����;q�"��ӌ�r՝� s�#�=����T�#�-�p�#8�"��%��v��!�`�(i3�p��ν(C�IחKD��ݚ�Н����(��x�Z��x�J�J�~>EX!�`�(i3KK�+��o�M���V��+��Q��:~����t�Ƥ�x.�Knq/�r�]/2�ݚ�Н��q�9�ͭ�M���V��+��Q��:~�'DV���b�z'hۉ)��d�7�q�!�`�(i3�����!�`�(i3���>]&���F�x��&���ő��̼��CH�+�e���;�z}+;��ݚ�Н�fĉ>99��j���Gp!�`�(i3@�c��F�x��&���ő��̼��]���J�"'��&އ��-/a8!�`�(i3�H�����kv޶Gl�e���;X�W>�V��ԜF��}�����Hٚ�-����!�`�(i3�'��o�u:��_x�H_��#���=��f�ae��0�U+�qbp@�!�`�(i3՝� s�#���k$ !�`�(i3|�au�(Z�H<�2�8��C"���h�G KH�F;p�	+��Q��:~�8w�B!�`�(i3$f��_Ub�F�S�1 �
�:qEp:䩒=]'!�`�(i3KK�+��o�M���V��+��Q��:~����t�Ƥ�x.�Knq/�r�]/2�ݚ�Н�����l��2l��*��Sr��3��ő��̼(�̖edЧ^{�jMdGN���!�`�(i3!�`�(i3+�&�B=�ޤs6Ed���i�4(��X�3��?-'��-����!�`�(i3!�`�(i3�5?�&P-ߑ������E�g�������(ӈ���m�r����!�`�(i3�/��@���-��(�Ļ4��aA�'J�A7���ݚ�Н�!�`�(i3��jVѭ@!�`�(i3!�`�(i3�5?�&P-ߑ������1��-P�͹9^l4zױ>������!�`�(i3.��J��__���Le��fi��W@����E�El~pDa�8w�B!�`�(i3fĉ>99��j���Gp!�`�(i3�	��x��ݚ�Н�!�`�(i3K�\7}�W,�����`��5?�&P-���ݵ����yM������^�|�3A�)Oqn�����ea��}Dq�f�!�`�(i3�5ߧE4��!�`�(i3�	��x��ݚ�Н��/��@����Tٷ��Ő����l��5?�&P-߷��Ѹ�f�R��ӟ-���[��l_!�`�(i3�5ߧE4��!�`�(i3��Ě���ž_�F�$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vx܇1~�}��Eg�N>Z�Cs`��)rʈֺ�/�X�G[��ht��R����A$�P������5d�	�+�&IiI9�o«IX0F�M���ѻ�����g^mb\���F�`yx�>�+X�[�G���K!�`�(i3!�`�(i3NL�Sfo�r��n�"��Wr���,(��9�e���}��G%�MP3�_~�:N���nF���<�W�.�P�	��
�Q�}i�]ʺ�
ǋ;�-mO�J�A7���|#HK���؇�M.9�[�2!
f������z�k��^�1��dc�@c�����h�'�ɳ��<�6�Q=��ž�Ć�T���7X���c�}�:
��x�{�\��N�Ś�-����;�jmT�#Q���V�_�mS8<�n�ݚ�Н��$�`V1���j;9ek�I����~uK7͍��|��W&":�ݚ�Н����F1��h��;��I����~u!�>!��!�`�(i3�����A_�͸ޫ�(��$�\%e��}Dq�f������!�`�(i3��ѯ���Z.Q�NJ�zQ!�`�(i3�H��c�L1���`��1tSjv�!�`�(i3�>�u��8f��P����'�^�����ݚ�Н��H����̲�2�!ڴ�4FF����w�FB��-/a8!�`�(i3-�E��%�w�=�J�5n��>�my$�N��o�/���;!�`�(i3��w�w:�!�`�(i3`
 ֢���@�k��}Ǒ�e}5���&u?�F���m¡!�`�(i3�5ߧE4��!�`�(i3�+��9,(�6� ;h$	�v��ONH!�`�(i3`
 ֢��.��� j�H]����j)����r^!�`�(i3h,ID��.2�6� ;h$	�W�L�sQ��|`��'��>�4N��[�1tSjv�!�`�(i3���F1��h��;���_r��Ӝ�}Dq�f�՝� s�#�h�����{"X��U)�D#������S�<Ԣ�7Z�:1�\mdЧ^{�j��-����!�`�(i3a3@��[/���fg�p5ϫ�X�>���8���&�
�:qEp�h?�4D�Ÿ���H�$��XCp=8�b(���sjߢiVr�r%)cA9��9dJ�!�`�(i3���Ȋ�?Ӗ	W��e��*}���C&��!�`�(i3�5ߧE4��!�`�(i3��Ě�����}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍ�A��XGX�W/��WuC=2崝�m�Wd�<�g�IL�E��6�o8:4�I���c�90�Ǘa��x���+�^n=\f�5>�+���B��d5%����aV�9�A(�c���_G��Hb�8�u?��I!�`�(i3�d���a؅q$��.��m�f.���G�?v��� �+��R�����ߠ����9
4�٩�I����~u���NM���A��4�h��T�?Z�k������8���[{/;k+Q�h'�Ȝx�5W ��̫(�8�u?��I���?B��#Ɵe�*|�÷�Wе ;�jmT�#��"����G��Hb� h�ҩΏ��^Kho�7�j�Γ��-����!�`�(i3�G����ic)�̩�?D�8���F{/�����,([�y�����ִ��}Dq�f�8Uf[���!�`�(i3*�˜	���.��� eoK�UuA�����5��x-#[x�I��״ڹ�	W��e5Z	�R/*__���Le�Z6����pK�9�b�u-/���y�8��C"��cG���`ö8�b(��@��C2K��NTP]�0@�m�W#�UK���6����>�4No)�T*�c�ı���X>��L��;+�'ն������|�Y[�Yy�l��A�.�� h�ҩ�
�:qEp0���Y$��D9��ɰ���|e"�Ra])n#���r����}�;��������/s9��$�\%e��}Dq�f�HN��R��bP�63Z�t;�jmT�#��|>��KK���������E�El~pDam�������ݚ�Н��*������Э~���V'�^�����ݚ�Н���w�w:�!�`�(i3Ɏ�#���?\a��4�%��v��!�`�(i3��Ě�����}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍ�0Hl��?��B�бuf9����� ��PdGZ鎬�������(���_C�/b# @�k�EE
��$C�~x���yM�B(p`D҉̖�7�j2��,zc��Ŕ��T�\ ��z
%3(�Z���L��O��l7������3m,�$�f^��h%O6]9���tk�Oȑ���Rl�Vn
*����!�_b�ȅH*�#Rn��'��9�������+M���<:� �����"?��A$�P������5d�	�+�&IiI9�o«IX0F�M��<:� �Ͷ�2��ibs��2[�a��o���zM#��m�!�`�(i3��4h�=Iz~r��V�n��dK�����fF0��q�\E��0�c.��V/ ���we��0�U+�qbp@��߆�p�h��d��JXl'�T��~��?u��C@!�`�(i3.�
9� ���(ٗ.;���JTv�䵶
�t��T&��ۥ`�M?��y�!�`�(i3�!AaiT��G��Hb� h�ҩ�?V��j�c�_�Sc��E�g�������(ӈ���m�r����Ra])n#���r�����+��9,({~1JS�K{�Kk	|���e��Y�	9צurT��-����!�`�(i32W���R0R�8�C�w~�h�8Vb5�!�`�(i3�5j��`q��+hX~G��Hb� h�ҩ��wӨj]h�H\e1E��v{��lw	޸���P7�ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vx���Db^���V�~�&�pɒu����(��gb#�o��_�Rv�䩲$���dS@Ɵ�o{y����i�q,?5q��7���9�hm�ko@h�r$ɓǃl[�Ƶ��I�q����!�`�(i3�� л�4�>������9�@f���ʦ�/\<���tݻ��=����t��p��b��_���&#ݟJ�a$�Y dN�<@Iv��nt=:��:5A��p�#}�{��8y�R�VN�c뵣�E�g�������(ӈ���m�r����b~y� �z�q�5y�!�`�(i3k������8���[{/;k+Q�h'�Ȝx�5W ��̫(�8�u?��I���?B��#Ɵe�*|�÷�Wе ;�jmT�#��"����G��Hb� h�ҩΏ��^Kho�7�j�Γ��-����!�`�(i3�kv޶GlWw3i�|�/ ���we��0�U+�qbp@�!�`�(i3��=m緒rQ����u:�uݎ0�{_8�Y��=�}�Vݨ��}Dq�f��� ���m�HT�AY!�`�(i3%��v��!�`�(i31���~�B�'��a���p��b��_���&#ݟ������ҭu:��_xV�PL[���ݚ�Н����(��x�Z��x������&G!�`�(i3|�au�(Z�!��w���N)_�7Z鎬�������(���NTP]�0@�m�W#�'�cL3��ݚ�Н�$f��_Ub�F�S�1 ���0���>����jP4J�!�`�(i3�\\�a���QF�����$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vx���Db^3��h�]Œ�i�hO��J�a$�Y ״$(�>g�����V���I����~up�@OM.Ir��ݟ��Da \6��.���v� 8��l[�Ƶ�%m�Y$� 1�#*���C5K�@�/̷_��yC��S8��4�J	~�p�����5?�&P-߇Vw��o�'���Xw�j�7���5?�&P-�O<�aZ0%�FQ��ݢ�^3DAf2t���a lI���;E�@�� ��r��x�l��1:�N�*�x�6�5�p���PF��W�!�`�(i3!�`�(i3-��<�ξ�\zǣ©��qr�^*4y-��u)+�*\��Mh�!�`�(i3���K�7���[�쮃���=����t��cg3/F�C����:�,x�~!�`�(i3�b[�u2�Gp��bە��Y��j3��� Q�N��*�������)�ak�m6!�`�(i3,��O^�{	��O� m5�s�٩���I��������|�!�`�(i3-��qW8+���ǣ©���L�K��%<7�`+Al��R��!�`�(i3���K�7��,+$\�M��Ỷ �U�
.�Ūz�/>�"�Ax!�`�(i3!�`�(i3-��EfVNNaJ �!,�<�W�.�	*}���!�`�(i3!�`�(i3-���i�4(��i缔]����=�<���XΚ��!�`�(i3!�`�(i3!�`�(i3X�PC!`�|��K�z�&�C�/��b�-W��^[�΍�>!�`�(i3!�`�(i3���K�7��+U���m_Esw�E��Wʁ���p�B�E�!�`�(i3!�`�(i3�X;p`��;���g��f�?ǉ�=�.��Ԕ^�|n�M�!�`�(i3!�`�(i3J�]�RU�`���,\ͨ܉p������aUMf�n�Q]�����	!�`�(i3�����[h��f\k`�k	���\�I�\�,�Xʚ@h!�`�(i3-��<�ξ�\zǣ©����>\�${lZlX�l��)��40� \��M��緾7�� ���&l@��8���_�[h�q��d[dͤ���!�`�(i3!�`�(i3�X;p`�p�
9��x`�|��K�z�&�C�/����o��,�Xʚ@h!�`�(i3!�`�(i3;o���D�@��;���\��f�?ǉ�=�1�)�c��!�`�(i3!�`�(i3!�`�(i3�u~xgA���������6%�a��<H���B�r��!�`�(i3!�`�(i3�X;p`�ct�:��RE3z%�u�܆����>[Hs�?����H�Ud���7!�`�(i3�&8�,��X��N�'��ҀL���G���ȍry��	� 䉇o�M���w0�!�`�(i3!�`�(i3�[K++�2�^����&Z>0�!�`�(i3!�`�(i3!�`�(i3�X;p`�)R��L-��竷b��"&�ڶ|e��!�`�(i3!�`�(i3!�`�(i3�˺�Q���f�?ǉ�=�-���k\�!�`�(i3!�`�(i3!�`�(i3Tl�������l6��'�al��p)�ak�m6!�`�(i3!�`�(i3��oC���:��j�g��Qc�:I�J�a3mPy�x�6�
X!�`�(i3!�`�(i3�X;p`��5?�&P-���Bx��mK�#]2��B�r��!�`�(i3!�`�(i3-�������?V��j�c�Ud���7!�`�(i3!�`�(i3!�`�(i37�_M��f�?ǉ�=�%]�N��!�`�(i3!�`�(i3!�`�(i3�����J}�b�Ot�i0�	�:]Ip�8Q"y,3@97�����Ѻ'�,�9�{/N2~-ٲ�5��X��?������U �Y4�@	�u�a�)���Ir@���Ɉ� ֒\���{���Mn�l��5�9��J�x����>�=�孒Е.|���.ն6�φ��<�6�@a� ��fFMqlg{y����i�q,?5q&kT҉­���Wl˦'ž1�|�'������C�ˤk���c0zQu��e��OA J�3���y�my$�N��o�/���;Sd��Pt,��X{2���q9+t�}�@��v{�G��|<:��;�P�8���[{/;k+Q�h'�Ȝx�5W ��̫(� h�ҩ�:
��x�{�\��N�Ś�-�������vo�q"���y�(�R̱�A�0���q"���y�QF��������jSA�q$��7w#NݬKomy6l6����|<:� .v+�;�jmT�#�UMg�chb~*��s�:;P���{~1JS�K{&�U��f����Fz����c0zQu��e��OA ��jq.k�e�kp
�:qEp�;�P�t�5fĉ>99��A0ok�����F��O�\E�W��4b-Ukc��R��4AL��΋I~m��D�Aa�R�