��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lV�t�[;�Z��4d���Ġ���딣0&_���X0���2|	p��rw@	@us���t�]�D�"�q��yq�`݊�|���"rG�
���}�\���V�S/+��K��������طǪvWa.�U4�,3���\.�"�K����u����l�|���j�I�?g�f�;K�y��rk�gH��(�_�|��2Ee�Y�R2
�I.��	���
���s}��=M���c���X6(!2��탯;\߰����G�;�r��1
�#����K�����MGD1�/��	m�Rn���L=`=ű?�y��D.�1o��������X��|gߦ^�y�b�5�!�� %	��}�Mx��+gb�Y�>�E��J�}�aE�d��n�NQa"_��ګ��E4_N*D$H_���HN�ۄ	B��]�A��o����j�� �X�����Hu���M~IMn�Bɍ[[B�����]a�{گ|A�U�O��g�k�q�M�4��t��d����G� �NUD60L�8yI���(	_dxd�%�GY�i�[��OI�9g��گÉ��`��Cm{39��ꎸ�W�����選��Ъ"�\�%�Kw	�Fҍ���D1�m �n�<�L�k��\"�!ҝ�U��'���K�dS��N5���oKגv����n�#��iM�j+�TM`�O�C��u��
�?�6�2��fs)�S�	s������0��+ȭ
�%��g0���CxU"i� [�W�a��X��١:� VrV�]qwR�	St�{�Pt�yhY4�!�����3�5Ὲ��7R��+�+5�:I���f%%eZ��T��B���d1���qp<}P�]�2��ӿ�3����óQH���1�@�?r��\�j�s@��:�����:�q��>p�.�o[�;ιV�&��'$�*�
����%��d�mVe����ʠ̴�X�S{D����ӀS�Ǩ�,�g�E��f.���*��ƣWB3��ub %���܏���� >sX��f�o*%�\h0fjˌk_ڍSSt�+E �ؖgP��c{���(���sa�MI��}Vj̔[�u�(�`��G!�W�����ħSq����@�����S.1������b0�[X�b\g�=�7�B�����N-�_�ӏf8�r\<%|��T

�F���W�� �D�ߏ�M��I�bI�xS"PZ}J}��`�{���GO���6�;�fy�F���F�bAg�
d�mFmDj��~�̤뢲�
29�/SM.P{�p��=7v��욓��źy��Ld_���"�ٓC�KI[29Tf660�(5�DX;7����A8v�[�L�9�;�7p=J�Z�Q7�=�'�*\޻��W���)��	3sXRC���<<��I\2�}��s���{|K��h�����a���5�FF� t�e�=�ݭ0���CxU"7��Y��d����) �o!�`�(i3�B��c/r��T��$.��H)q0����K�#B��?^
ر��ZXty���`�c�~e�0�We���ܮ�c:��1��q������-i����^!`w�� ��A�]�B=>_�o&�8��/M4#>Y��<<�٤:�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��r�����A�F�7���3�GXS����E@��~���($�J.���
�=W�֯��i@F�5�=h�GD����c���o�����0���S�BgV�0�ם�k���s����Ct�z&��ÃlO ܅doGa�젿��ʐx�?WA{I�Z�T�����N\� n��A�T�g�v�;�K7���'n�^0o�)�?�^�?�XW������w
��ڎ:�ڛ)
�}��ɣ�YV�PD�E${��4`�˨�;O8�d�
~�n�}Y�:]�@�<g��ũ,+$\�M��lJY�Pt���`��8��f�`��[��Yt��'�d"[~6����aD6&>��Y��q��f�}��`<Y��sp�����5	���]���c�A�L'�������W��_�ړ8���/��4��}�<�N컽kg����|g�Y�'���Xw�j�7����'�e���"j���b7|#9���\I�d#�(Iѧ���i`�ҋX����>��l%i�-�M�g����Y%T��BPe.��xu	�>��l%i�-��9��稕Y%T��BPe.��xu	�>��l%i�-̇i�d�?�Y%T��BPe.��xu	�>��l%i�-D�wP�/�wM�Ǿhm��@IE�U����S8�
T�F���u�܎����k/��m#�U��_D��.V&��B֥�(����5��M�=��S�\��3t��Q�L��w� Oag���:tӫ�C+��T���.��Б����K��!�9tf<[
iEE�G+�T�J��h�H�MPq6.�b9�����6�_��1�m��'A>/y,�Z���rS�b�8Z���'�e�����"�?;(��j67�=t�!��&r���q� N��p����IÙ=�Hʆ�In��t/p���xL��fl���=��fLR=t�!��&r���q� N��3�AŠ�zL͊�q��٘�27!�g?_��<'P��!jcCA�T�g�v����fQf��p�m~|��4FV�{E�JHn��z�'8^�#ٸ�U��֜��3Ԓ��������\6��.�E�]��c8?-+eN�s(^��^p��nk�Y�P	dU�1�1�����1#��Z�����XP�����'�e�����T�LJ�n��f�e��}�
�?�`<Y��sp+N�f�+�n`5�fK��0z�cUL�?m ��0���k��$a(􆿳���2����.��DP֞ �T�'Y���A�? ��p�]�!��	Ǹ�y85�����S��Cƃ
ᾆ�x�T�\ ��i3�|)sՀ�T:���V�Z7����6	зq8�Ј'���Xw�j�7��Po�Q�>°������R�wX��}�
�?����2jɸ4�r�@E�n`5�fK��0z�cULn�4Z_U���l�����"X��[��Q[R�7�����bpZ��	�`DÜk�K��h�d�٣��c�A�L'�"��/f~�\	��K(����`y����@����gG�������E3-	����#�6�3��rs�i�_n����B�Pcsù��Q��Y����2����..W���ۗ���WYHpYyI|*����]�!��	Ǹ�y85�����S��C\	��K(����`y����.�����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��U(a��,n��#Y��0!!�?��-�(�r���K�������D"�Ե��>���G�Q���Q�s-`��|��f�&R�߷�C��x��;����s�{uN��;^��ooRm�J��@h�1��R�������
��J��9�r4 II"��'N�����d�x.s�2��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �L5ӥ����2�l�\��#�ڊ<?@���hWG�K� X��V엽ߚ��u����WYHp �:�Z��pb!��u�^��po�����A����|�������-�YM*b��93�|q��-��kѶ���� >�������d
z����YUr�(��z�j���l��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ���?-n���2z�W0i��G2'�{�*��<$[S���=3݇F1�k2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc0l�f�m��џ�1�?"�MC@���U��S����k��$a(􆿳�eJ�Í6�UW��7(�bO���e�[i���⬮1�����ׂ�⾉�ƃ
ᾆ�x�S�v�b�k�#7ۏs|�-ذb�F�x뛀��⎽�?kg�w��CF��^�ߨ�,R���"X��[��Q[R�7�!#��Rh�1_!��Xm�`�V�s�p��;1�˚z����'6���;8=�g��U-�ePo�Q�>��	�Y2�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �LC�x&�8��*�&�.�w	�G�ԋ׺@��ϓ�9g$v.5�,^��o�ѽ��L��[�1��4��}b2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �!�P{� f.�Э]&k@C�Ɨ0z�cUL��ddՅ<Ta��;���=�[%�('T����7 �>5���P�ڈ�KK?B�5 �8��B<�·� � �uw��o�Ķ
1'�F*�L��!�`�(i3!�`�(i3ouD�����rs�i� S�xSVeb6vJ�pZ�*
T���џ�1�?"�SҢ��+��*)�2�"ղ]�6��21SǸ�v��ZZ>�ڗ�\�����V�5YZ鎬�������(����.��$��Z�d-�~E�`�_�y�1�����b��[� p!-B=�6f�0��>�;!�`�(i3!�`�(i3!�`�(i3!�`�(i3X�o|3��b�Bϱ��!#��Rh�<Q�vn��l����I�/=k��%�W�%�Ko
�S2�	���3\�a�C����e'{w#/ B!�`�(i3!�`�(i3��]���c�A�L'�ɻ�L�1p/-��ս�9�j�����oD�d5z�R��5 �8��B	�PT����َm(5!�`�(i3!�`�(i3!�`�(i3!�`�(i3P"G�wk�Z�d-�~Ee�1���1�����b��[� p�!#��Rh�/T��o3����f�RE3-	����n?�C���Y�{'%s��$��S���b�Bϱ�!-B=�6f<Q�vn��l����I�/=k��T�'Y���u��9�!�`�(i3!�`�(i3!�`�(i3!�`�(i3h큈��]v1�_ُ%�W�%�KY��{&���'6���;8=� ��g�SE���̵?o���$�X!�`�(i3!�`�(i3!�`�(i3!�`�(i3� �
{�������'}a��	����F*�L��!�`�(i3!�`�(i3ouD�����rs�i� S�xSVe�W�6?��W��7(�bOpP�Fc�����k��$����导�?!6)X���M����N!�`�(i3!�`�(i3!�`�(i3!�`�(i36�&��=�'�)�Բck�A#�G=���%A������D�ϲ]�6��2g�1�9�U�)��5npg!�`�(i3!�`�(i3!�`�(i3!�`�(i3�<�0�]�`���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}ں��D�&�ߌe�X� G��v�u9�oݮC^eG=2V��Q�W��	]�	3Y��P4ozz_=�\}G+�m����tw�$��%*��o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cb�P�z���5|����t�T��?E-h��$^(?��"]�B���[:Fa�7��M�S�"���2�y��|JS��^�uJ#��r$ɓǃl[�Ƶ��I�q����!�`�(i3�� л�4�>������9�@f���ʦ�/\<���tݻt�{#	�x�_�Qf%u�n��>�my$�N��o�/���;�̢k���F�KD�Vr[/}>5��0�7<(�lb����y��lD�7m�T��Ʈ+ˀa��z��2�,�$XR�QܛOcOZail������&G����l�陜�f��D��&�%���>���@]�'����u��r���2��}��e�g��)$<��0n|�!h�b���t�lE�YK�f��i��#7ۏs|�L;Л��|#9���
�:qEp'{w#/ B�2��}��e�g��)$<��0n|�!h�b���t8L��e�x�f��i��#7ۏs|�L;Л��|#9���
�:qEp�;�P�t�5fĉ>99��A0ok�����F��O�\E�W��4bM�S�"���2�y��|JS>d���9 $)�lj�iE�EYZ/�.�L�����