��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��:%��Z���xN��g�.H�{�|�w8�M�Q�"�,�#ѷ���� �\_I+ĂiW,���D�+y[ف���rn��mo����/~.)��3�(����C�X��2�k(����)O��Ξ4�"�\�� ���K�O�{�������>�pÔ���c\֣�I��B���t��|U|�/֚W����͇M��Zw�U�;�\��^�� ���K�}M^UQ�S��)�e
�9��Ax!P����,��*�b؏�@�~�S�`\��Yi?��n;�|-���g]����g�����fP����IL�+��ץ9�^kh�u��<��T��� �}+~�8Ó B]�pE(���B��|/~.)��3�(����C�X��2�k(Qg�@zh�S҆�|n������}�K�~^T�ɴ��b��9J�Й�m�z\H�� 0��~����p�:�C��JS�Ȕ*Ĥf���J�D{g�P�r�|A�l&K[�
C�9���1� c��(�U����	x]�m�Je{q��P����>�]!�ՄN�Ӿ��)�$�����PГ��0�w&��EO�{�������E��sޜ��*�c�N!ͬ鏈wƠ��ѹ?�����qU�%��Sr�'hJ�.;��L�OT�+?3�l� c��(�U����	x]�<���e��8�t�~��,�O�W��s�!5�S��H���)��������ҥ{E�?HF��eUٻo���mi��*	�ť�.^�i��' 1wH�x�xs��3�<A��z����
a�������~�+��,/,����W >g1�]l�&Y��F}갨y�����# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��`y��f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�}�Z���ik2)�
}wʭU&H�1��8�h7H�u�ÍeRuw�C?3d,f$�7Q0�"<�F�ٴB�I�SbW�{b�2"���Bpш�#w��s8[Z�xZq��t�1�:�Ω�`<4}��o�r� ��J��ݪ�nP;���7	�\�Z�م�L�Xڈ*-��]���P��`�.�D���J7"H�f�J2uZoO�=���@$"��ea�8���*���g S�ĲW��,)�W*g;X����ˉ�1�:�Ω�յ�'�)xE���8����s����Ct�z&��ÃlO ܅d^�R@Κ�2X��9cѶ��[7�d|���XP���4֔ʽ�I7��-5��3�Q��\�vņ�Q�]��8��ؤƼm��P���ݪ���[7�d|���XP���<����k�|���0/ܤ�(g��V�[7�d|���XP���A�����L(\Ӧ�$�̎�)NC�lԇ�-{���|g�Y�'���Xw�f�VHF��Q�#<4^���|g�Y�'���Xw�E�i�m}6�B�r����|g�Y�'���Xw�4��}�<������Ə+k&v�Iz��j���'b�t	�U���C��O]r�<Uee��0�~?5+�&Ã�M�R�^Ƒ����"X��[��Q[R�7�� ߌ�ˑ����E��@IE�U����S8�(´W�w#�m��P���ݪ���CyW�f�t<|����faՊJ�e:[e��mea�8����:%��Z��vDY�όWU2_*ϝ���67�a��c���}��D���(��z�j�)�q��1�:�Ω�յ�'�)xE���8����s����(��]��'��wb�*ܑe�W����n�4�c_����+#��.X���*"v%)��Qcm h�]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e,%�0g���[�=�5x�� �i�#n����-�*ܑe�W����n�4�{lGD�V�B�9Cd���*�=��X�FP�=��p�m~|�֫Xaʬ�����]0�mt��e����#�wb�S��V��\����0u���g}eY�e��Hz�ay��0�~?5+g^�z$OO5b11��m��0�]cJȷW+`�x�o��7YI9�D�@�Y�4��j�O$� ʳ?��A�Ws#Cr����it	�TU����z~��6��	���`y�����g�,P�n����|!���^��\i�@^7&ģM�2�T�������it	�T���-M+�Ԍ���ͥ�#�><,v�;�@����gGkx[JaBS!�`�(i3�6'��-��oP��a�I�v��9��"�����BȀ�������Lr�u�Y�KG�ξ���X��9cѶ�E�����+T5�O�%E#P����o�af[��C��L�Q׭n������.'�'�)�Բc���W�g-�R%�����it	�TU����z~���D)9W ����,�ǰ��i��W�ot�KH��p���o�P٘Rly��;U���2�9S�Ɵ�7�OT�,���t�\~R�W�u%+�$�M5�O�%E#Po�|MI�yb�V.�[��	}�@����^Ao}��!�z�� !R��0j`����OD5�O�%E#Pd�G}%��Ď��J��QCT�"�x9�¿Y�����'�U$��Y�]5�Z�z�.��7]���boNF�<}��!�z�� !R��0j�^�̷ؠJ��:����SƏw0����QJ��-]'\gWg��	�Z�kfc��2���8[����㹭�o��7�!�`�(i3xjzӝ���I(͂��-����!�`�(i3����o�a{�C�/pkE�g�������(ӈ���m�r����
�:qEptiND�S���/9�=eSe.��a��o��ѵ��.�~<�Ɵe�*|�÷�Wе !�`�(i3�s�Yls��8��GM��-����!�`�(i3FkH��۰H�J�����Ŋ5�m�/)+?����$�59�
����OwV����Tׄ�~^�������v�ݚ�Н�fĉ>99��A0ok��
�:qEp�;�P�t�5
�:qEp$�)�vxk.Db[휯}Dq�f�����,�ǰ?%{B��0B�.��(�w!-㫓L�yF�=N��އ���$�d��4B�%iۋr(���w�Ε�(sہӛ�_��s�֙7�}�!��ނ�`��\y���t�T��?E-h��$^(?��"��K��O.C��WHe�Q!�`�(i3�'ž1�|�'����u��r��!�`�(i3L�^��*�d�:��5c�dN�<@Iv��nt=:��:5A��p�Ra])n#�璓�c�������t �[l;[�G���KlG%��`��ǚ��ظ
��@�U#!�`�(i3܌;���'����u��r��!�`�(i3����o�a{�C�/pk�� �X?�V�BHS�/��
4�e �S�!�`�(i3HN��R��bP�63Z�t���%>�rGO�D mWN���%>�rG߸��S�Ȍےú9(!��;b�-�2�V��	��y$���/`�K��rw.�g3Zv���� 5i�
�bx��.�g3Zv���� S;�d��3Tp�m����&k@C�Ɨ0z�cUL��Zi+�E�j1%vN���y���_gv*���h�b~��Z�[������H��<�C�Ar��� �9Cd���*�=��XƂf>x�:	�W+��W�A�~����Ձ�=�n�4��Ǳ߁R�^Ƒ�өwo��Z��Ac<�p{�5�O�%E#Pq�\E��0����E�I��#ɱ��<��>��𱒁�"ʥ}cG���I��)���W�w��fDU�����.��;_��8W�w��fD/��6"�^Rr������%�<�$