��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��k�	G���D7@aI|W�ϛ9�� ������[���a�8%`��4�s�6�XAoeuA�D3�O�þ�V��vMcr�|�zc`�G?q4%�}||�'�U��P&;m��Κ�P/�u����)O��Ξ4�"�'Y�L(�K�O�{�������>j� �`�c\֣�I��B���t��|U|�/֚��LT�E�9��h���$[Z�i��%A�a��gs|�e
�9��Ax!P����9SA����q�HS�b"L]$7!����Y�f��a�Z��Vׇӭ��!�`�(i3h��8�|�g"#~j[O\ڀB��+ H!�`�(i3!�`�(i3�f��)<t>���PF�!�`�(i3A�"̙��2�����Vc2�����Vc.|�('��r�dZ��߉�󆭋;2�����VcЁ=�t�!�`�(i3CS�Y%��t[Ed�+֚L��2�����Vc2�����VcϔJCS��G�d<��2�����VcpNR���b,�ҧ�ɟ"Y|fN�:@��翛Sf�\�_�Ճ܇���'o�fqII��*�T�٥��T��|g�S� -E�7*����q��jlw��JF#�dnE��k~xhd����Cr��1��i�Vw�oM �%���bv.�]ֶO�4D6=���i��p�b�G!��Z%�6�ǀg��i��vp�\��M��ڀK�_�rۈX饿��!��o���ݯ_gWgj"���\r��3ة�K�~�'o����֜,ӘkR� �KF
������:��ۜ������;�Ӏ��B[/'g�`	�K4̓������9(���'�Pw��[#M��*�v}���<�LK���i�[-z�g��hs��%�-h���C}�{�c\dnE��k~xnE�HC+��3K�<�s�������5��w�:j�.Ѵ�����T�'�"�ݥQ����2O��'HY-(�3�(M���O|x�Ͱ��Y$��7\F���r��RL�a))�kc�߇���G�/9'�$���'�r{V.� !�zg�Z�$充�pje;��M͝75#S9��%V��"����ʉr���u��w)�Sl���-�ed�~篟|��d���Y��^"� �/Jџ�_�v%�����:��/�|^��D"���b!��k�8���҆�|n����wH�L��Rl[���.���M�ѕ�����aWfL1�Q�j+�B]g������Ⲕ�u��w)�S�3k:�(�-X�7�j���,Ud8J��$�ƶ��Ÿ?%�b8�<�#�1-@��%��Ձ�k�8���҆�|n���)kd&Z0�i&��a�&����?ʳ�W�%"4����*�T������|�OA�
܊��?Y2���3m�!=�y����h�}D�8����8Y�&�\�#�W��a�erp����N�u���u��Uy�PD4KU7B�����<�[0YY���\�4�sP	�b\qB8Y�&�\�@N��B@��2�o n;�q�m���mi=��B�-x=�WD���4B'���S�K��i|ٓ������v9{�$W
?%x�+�� fג�� y�dH�]��/�2�-�]?�B�nI�4q�Qt!��c��<%>ì�oJ5�%,�k�W��T�٥��T�Sҥ��|E�EYZ/� c��(�U����	x]�<���e��8�t��s*ո{�x�G�F�����OwꅂF�-!d6߿��b��'�� |X��M��"�D�u���lٽ�G��k�8���҆�|n����{y�ڋ�jV%[&��\�۱��ѕ���Z�[�0�7٢z|Mߘ����g�/@�G��P�?^
ر��ZXty���`�c�~e�0�We���ܮ�c:��1��q������-i����^!`w�� ��A�]�B=>_�o&�8��/M4#>Y��<<�٤:�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��r�����A�F�7���3�GXS����E@��~���($�J.���
�=W�֯��i@F�5�=h�GD�#�̔"v��ƒ)?˳R����.��ѬL�1m��+Y#_WӢۉ���2=�l�����뙇�� E�ئS��.V&��B֥/~.)��3\�R�F*}�c}��uO�Go@3w�^�����������,\ަ�It�ఙr<	6֚N�<�x�]�V���&;]"�f���3�2T�c�$��b9���1��]2�?V�Ľ�߉��ə��Q�^�y�zL͊�q��UG�s���q����E©�ʐx�?�'n�^0o�!���!��6�e�:r�"(?�M�_뎱�:L��ҭ�Y�����[�����cJi��2�S�ڬ��M����@qzL͊�q��~���r'�+0�l�R<�q��f�}��h�'f R!�`�(i3c��Et��q���U�ЂDa��(o��0��7�����5	���]���>����C�n��J�
��Y%T��BPe.��xu	���S8��<�J�QM����2�E~9���i�d�g��U-�e�,���6+�{���"�,�>E����-��%Mό���.�س���*G�`�B7d�N�By3��<�]�!����M[��Ǣ.g"UƄ3�|\�x�Z��-��%Mό���.��D������A����N�By3��<�]�!����M[��Ǣ[��l�,�Cc�70�TD��ό���.Ӂ��̰�!�Xy|�WN�By3��<�]�!����M[��Ǣշ�G!�C"�,�>E����-��%M�rs�i�jf� l��E�4.@�7��y%%��`y�����:�Uw�j:��e+������5	���]���>����C�@�,{n8_�_~�:N�c��Et�Y�{'%s�ui�铨g��U-�e�,���6+�7�UyR�j7��h��;	�TD���rs�i���Ӧ�am�T�\ ��̭5i��2l�~�+yp�l�E����F7G#+��\w��0]R���5`j�`�B7dԘ]2�y�Z鎬����[�Rs&�ggy�т6�-��E����F7G#+��\w��0]�V�qZ%	u.$����]2�y�Z鎬�������(���pl!�6���;b��g��U-�e�,���6+��>1J���"�,�>E���TD���rs�i���`�M�	=̞��>����� +'������݃�Q[R�7�{d��L�>PiM �H��]SBÀc�ȉ����;WNCD?WS����}�Cb�WA|[�7��V-�}�߰S�j���-�7x��
��������E��@IE�U��>��l%i�-;�ƽ�/���AS������
L'���Xw��e��c<��7�L���5�N���p�@IE�U����S8�<�)��'��*�S#^�V]��}<|������N�?�_uM��y��I�+��T���jB�Fg�Y씤`��p}RQaI+k�U��OV�\���G}q�P ڨ��S���Qߵs<��7�m��+�<4��ˌ�ň��h���T�%�/ң��Z���y�뵵�
�$��Xo����HcTz�Uhw����\�v��\aьIR=���2�E~9���i�duKr�'i��g�,P�n�r��A�, ls��+���K�LD�K�T� $��We���M���!ؒGb!��u�D��ɍ�٠�и�0�G�w�^>��p3�+��m\���_j���5z����k[���g�v�b!��uፏ����V?ː���T[�Z鎬�������(���pl!�6���;b��g��U-�e,%�0g���z���Q���j���2˯�s�N��ό���.�}�
�?�ﺌ�<$2^��R#��]�!��11<�InN�0���ɵ2���HF3�@����gG��������`M��
Z鎬������_�,��LE-L [�/��$ʖT�d�٣���N N�S�+w�7�XB���2#�n`5�fK�\w��0]b!��uፕÀ����yPl?.���cY�~�"���ʷ������<\)۟���4�%;ך��C�:�S��0: ��q��MR�ۘY�{'%sAX���	q�KS���K����)��T�\ ��i3�|)sՀ��R�A0^L�H�߳Mkзq8�Ј'���Xw���,D�C�:�S����"c%�B7s�9���o��S8��<�J�QM����2�E~9���i�d�g��U-�e,%�0g���{.[��(��Y�b�΀�e��Ek�Z鎬����t��LJ��{�� ��8D�N������Q]� _�rs�i���`�M�	=̞��>����� +'������݃�Q[R�7}ϼ 8�������qJt� n���]�!����w�Հ�	�-�_Y��r-�T��v�z��]'���Xw�j�7���S�ڬ��M���q�tt�g��U-�e,%�0g�����9וP�;6�2�)r����'���XwI����"�d���m�0: ��q�"�k� ��Y�{'%sAX���	q�KS���K����)��T�\ ��i3�|)sՀO'�[m%#n���R�7s�9���o��S8��<�J�QM����2�E~9���i�d�g��U-�e,%�0g���z���Q����by��Fзq8�Ј'���Xw�h\K�5~�Wv�A��2���HF3}�
�?�/$�ߺ��]y�ei��nZ鎬������_�,�;�7���c�eK�	�$V�7s�9���o�jƓ�[b!��u�lv0�9l7s�9���o�jƓ�[��ǐF��nrm؊(��@����gG�*J�K:�*g�YӅ:�7s�9���o>��l%i�-����힅	]Q:h�E����FZ鎬������_�,�;�7���c���=�ڹ&��Q]� _�rs�i���Ӧ�am�T�\ ��i3�|)sՀe)����|�>Ht�u�U��Q]� _ό���.�}�
�?�`&c�'N�j��2Dg���d�٣���N N�S�dg�W�p᢯��0�f��"��'���Xw���,D)SX�:�_�o�@^0�W9a!@\w��0]b!��u�ì�u"4�"�,�>E����\�v�g�W�I吱 �']g����
�2(�;���,DD�=�G^�qe���b�l0��F��jBo�A;h�F#"�G���T�c�$��Ne;�*��9W������\�+�J���q���U��@����gG�	�L���0Ox�%7s�9���o>��l%i�-5�e`��9G$�ء��E����FZ鎬������&.*O_uqcW�(u�" Oag�֠$b#^M�Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�ˊt��q���1U��3{@�02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc6^-Yu�%�n��UM>8c<�@�ׅHK�b�"�?�a~[�B�׾ŞWsuz֯���,���ζݧ��~�+yp�l����;q���N4�j�ā��u;s�e�$X,�;ޱ�H��z%�֕SM!{yR�D��Ø
�`o!�k�}2�0���z��[����{y�mV8��/��Q�D�T1�8K��4����U̓���m�(0: ��q�\0�W�$�;�cM���/Ύ�T�L��/Z�o��>��Z{��0����3�soL�($�Q�rV�Fg�YӅ:�ht��p���=�?�Ҹ^���S&�r!�`�(i3���$=����I�����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�%A#�@�N�to��h�T� #�3Ł1�q�7��N�6�Q�3u&����J�f���-����R��ݪG�B�	z�M���S�-I�!A(�"#~j[O\�&�����1�sI�Y����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�
t�������t�T��?E-h��$^(?��"]�B���[�.��|ȃ�A(�c���_G��Hb� h�ҩ�q�� �`>��s��k��^�1��dc�@c�����h��-����'�)�����(9�ϦZ�Be�A�}�	76�&�� Ӗ�t$�)�vx��۽`�$�l,.l&�7s5kL�s�)];I��K�&�a���3Dr+�4���	+��g��=R���>��骾&�2�0���w��_>d�����r�����m:{�!�`�(i3!�`�(i3��!\�'°����ԬQ����lwE��$5���lJ1��j�p�B䁒_[�Ff�?ǉ�=!�`�(i3�#�-�p�m
�ܲ�#���n4s1�U��B��-�ܜr�a���DQ�^�鄃��;��ʁ���MյV~LvA!�`�(i3��w�`L�P�~�9��}Dq�f�}I�6���N�Cٺ��G��Hb� h�ҩ��H����D3w��'��b~*��s�l\�=�]y��d��-��!�"ǉ�t�����J�ϝ�5�v�z�7s5kL�<��r�ŁH�RtV�^CH$�I��*�M/*�3� ���!�`�(i3��\ Nh�gdq�_x�ֺq٫[_�mS8<�n�ݚ�Н��� л�VZ�ڋ���Y�َǤQ�Ї�!�`�(i31���~!�`�(i3����-Jg8�iT��*��C�Y�\�fĉ>99��A0ok�Ra])n#����,����0�|��';��#j�ݚ�Н�VZ�ڋ���Y���GiL�~�fĉ>99��j���GpG�&ց�*�7�|�9��n�7�Y���_j������
C�ݚ�Н��K�,ǆ�`�íN=]a��o���H�RtV�^�Jo���jk���%�8�Va�ir{��b�b�*#o�]�ʄ�v�4�?zm�jd7}�� ��M�sv��>���F*a��o���H�RtV�^CH$�I��*�M/*�3� ���!�`�(i3�k��^�1lv0�9l�'����u��r��!�`�(i3��w�`L���ǚ����}Dq�f��߆�p�h�Cd��9s��'}����=��-����!�`�(i3�FW�DVx>74/���RZ�Z]�+����%>�rGO�D mWN՝� s�#�=�U�u�íN=]8k��.ͥ�H�RtV�^pT/�GS�7s5kL������� h�ҩ�9��n�7�Y���_j�����9�x�\M�ݚ�Н��̢k��� :b/�Ti'ƃ�3�Y1tSjv�!�`�(i3����-Jg8�iT��*>������fĉ>99��A0ok��fĉ>99��j���GpG�&ց�*�m*H�	9��n�7�Y���_j����I�����&�ݚ�Н��K�,ǆ�`�íN=]a��o���H�RtV�^�Jo���jk���%�8�Va�ir{��b�b�*#o�]�ʄ�v�4�?zm�jd7}�� ��M�sv��>���F*a��o���H�RtV�^CH$�I��*�M/*�3� ���!�`�(i3�k��^�1lv0�9l�'����u��r��!�`�(i3N�-�}q�j�֎����-����!�`�(i3�B&�G���M/*�3��GH�E<5�!�`�(i3CH$�I��*�M/*�3� ���!�`�(i3�	��x��ݚ�Н�9��n�7�Y���_j������
C�ݚ�Н�fĉ>99��A0ok��
�:qEp�;�P�t�5
�:qEpj�E}4ظ�N�Cٺ��������� h�ҩ��H����lv0�9l�'����u��r��!�`�(i3��w�`L�ķ@���k>��}Dq�f�HN��R��bP�63Z�tHN��R��F F�E̠(*�O�q�)����CH$�I��*�M/*�3��GH�E<5�!�`�(i3����,����0�|�_�mS8<�n�ݚ�Н�-��)'�>���F*a��o���H�RtV�^CH$�I��*�M/*�3��q�t	<!�`�(i3��\ Nh'{w#/ B!�`�(i3��S����=����h�[� �c��!�`�(i3��Ě�����}Dq�f��k��^�1���+1��*Hx�g���-����!�`�(i3Y�5�n�����_�������&G!�`�(i3VZ�ڋ���Y���GiL�~�
�:qEp�;�P�t�5
�:qEp�;�P�t�5���aR��ݓ�W���{��s�J��ݚ�Н�����-Jg8�iT��*���a���݄�倮(���������d9=���u��r��;�jmT�#�0M�Ŷ�Eʨ�`N/������&G!�`�(i3-��)'�>���F*a��o���H�RtV�^!�`�(i3��w�`L�P�~�9��}Dq�f�՝� s�#t��ۻz�˾ �����]&�U��f�!�`�(i3<�6�Q=�hNNR!���	�-�ud��X縤�q
˾�'v����UrSuͫh�<���D��ܒT���.�[M���r����!�`�(i3�(�d���Հ�ˤ�䁔�`i�����tZ>P��]�{iK���	����;� �GE@��!�`�(i3VZ�ڋ���Y��ˇ*�h��!�`�(i3���F��O��ݚ�Н��̢k����0M�Ŷ斗���%�������&G!�`�(i33~��d�Mkٴ�$a�DkW�����JӉ��;4e!�`�(i3���ܚ��@��f�\%�~��\��8!�`�(i3�5ߧE4��!�`�(i3�5ߧE4��!�`�(i3/�"����V(pyL0DMlE'�! CH$�I��*�M/*�3��7ݽ��!�`�(i3}�	76�&�|��3��׹��ܜr�a1r8���I����ht��ܜ�[�^���H> �D�9�{*�,6����Z9��J����*��m4�b �	H!
�I�N��M6f��,�,&�J�����7�y��ħ���n��$z.��X� 2!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i33��0�����+1�;�.��1���,:&�����9�Ԇ��|Z�.!�`�(i3!�`�(i3v4{����U�ɶ)Z�_v(��ڥ����Ⱦ��,Յ�1���~!�`�(i3?Q�@X>#�-aw�n�W�^�|��p�@OM.Ir�H����2��b�Bϱ��>1J���� ��0� 1���~!�`�(i3?Q�@X>#�""Q���S=�r?z�3� �mKgN�쁘o	�V�6�J�J KB�~�.$d�I�vNR[��j��d��\\N�2߄��`c�N엁�7���R��4�{$�^&��AՉ������b�Y>�fWj�t�[LY�ЈɄu����0��|͖Dzd�=�/�t��Ǽ�d%���P�.�5k��~��/6�o8:4�I���c�90�Ǘa��x���8-|�D���"sS<�0�zG�������&G'9�и��{4hz�<Ρa�E�Rq���my$�N��o�/���;�߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#&�|Ξ쭧S{#�lܵ�p���S��íN=]n�|�-3�lv0�9l���ў�L��X� 2���t��Һ'��b�%���!j�l��XulMd�[���}��M�?L}�7x{^4��*m!�`�(i3�����V?��	����pॻ}����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍٽt� $�N�����"���Q�������t�T��?E-h��$^(?��"]�B���[�.��|ȃ�A(�c���_G��Hb� h�ҩ��W�3�-6�n��j&b�z'hۉ)��d�7�q��k��^�1��dc�@c�����h��-�����Zj���
���+1�;�.��1��!*��*8��!�qg�L�[\�"��-����;�jmT�#�[�#��w� ��Ք��ݚ�Н�U��p��PrΌ^pG2��$�)�vx�;�U4�IgWaU �IH�RtV�^>�Q�c6�J�
�Mɏ����V?��Ht�!
�:qEp'{w#/ B�d�tuљ�FdG@/X��-�����+Ut���$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vx�qb�V�_2��Z���}��C˥�ɗ�iL�G��IX0F�MV�ҁGG%4vkz����`���φ��<�6����N4�,�7����r$ɓǃl[�Ƶ�1tSjv��[�	���d�~{��)P<�ܓ�Y�̢k���F�KD�Vr[/}>5��0�B� �b���]���`T����+1�;�.��1�](g���������lҡ"#�k�d�8��k�SA/��M����,�,&�����ᇱ�@�=%��d��-��!g��J�s��z�
1���;#o�]�ʄ�v�4�?zm�L�[\�"s)l໶�,3��0���3i��U��N��M6f��,�,&��$��!'Q5/�dI{��XW���!�`�(i3+��Fe���5��o*4�"ǉ�t�0/0`9N1&�2����1tSjv���������5)��Z^�h��N�M�ob�H���T�ì��������R3Y@T���אQ�B�<}׼����!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3U`�Ȝ�W�iy��*)ci���{2�k��^�1�3i��U��8����q �H�%��ZtV1{,�m���B� �b�Ћ����$�~�+yp�l���d�L������.��U)�~[��Q,��:5A��p��jVѭ@�mJ�0�6������$�~�+yp�l�#QSU:�����|e"���F��O�}�	76�&�� Ӗ�t$�)�vx�+	=H�ลGH!aߗ��.�����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���
�x^�LRXN+EWE� �����D���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcZ�)���,I�$�*�����t�T��?E-h��`f���sd�G}%����3f۪�G�Q���x�\���F�`yx�>�+X�M?��yЕd�tuѽ3y��s��>H�,b�z'hۉ)��d�7�q��k��^�1��dc�@c�����h��-����>�Q�c6��=�ڹ&��nF���<�W�.�P�	��
�Q�}Ql4�u��;	ȕ?�'����u��r��>�Q�c6��=�ڹ&XC�K�7(��gY6!�K������B�̢k���`&c�'N�jLm�<o��M?��y�!�`�(i37�UyR�j����^7��œсW��e�p�x��;b�-�2��|$*g!<�A�IS��03�� <I�����&G�����$ZtgQ�9OZ�s:�8��z�Ȓ��\:9�C�s�4���%>�rG�@�	����$f��_Ub���uQL+��φ��<�6�l�x8��-a=F�!#�&��>�quA0�e]'\gWg��	�Z�kfc�_	�Ƽ��S�J\70C.�>��V�m^݆��xjzӝ���I(͂��-����J>zߋ��>ַ�����ƍ2���l�����g�Z��3��a���!@�f")u��r��}I�6���N�Cٺ��#o�]�ʄ��.�L��w)��
=b~*��s��m���>G��Hb� h�ҩΞ �@[������4Yz����|e"���F��O��|#HK�� ��5%q���f�e�x��w����֯���,mk��L��a�	�Z���ވ��*I���b�Bϱ��>1J���� ��0� 1tSjv��l�de����O|���/��kOT$f��_Ub��7��G_���;�P�t�5�׹���8�2W6�[�6���"����)W[�ۺ�E�`�4�l�T�܆rl���CLmk����������B�s�Uo����~c��0���IX0F�MV�ҁGG%4vkz����`���φ��<�6�`&c�'N�j��v�����r$ɓǃl[�Ƶ�1tSjv�œ&|�9�n��~��4�)P<�ܓ�Y�̢k���F�KD�Vr[/}>5��0�B� �b�Ѐ�(���0���;	ȕ?�q9+t�}�|#HK�� ��5%q���f�e�!\���k���%�8�gVdxQ,#�%+V��t�v��ONH!�`�(i3s�Uo���ַ������?D�8����Ě����E�i�m}6O�D mWN��ܐ�}ĚȜ��Y���ۉ��K�A�a�ܥ��(J]֞��_�TYh�p��_����3Y����P-r�uh����s�Uo���P�<�^�s�IX0F�MV�ҁGG%4vkz����`���φ��<�6�`&c�'N�j8D�r^�Hd���"sS<�0�zG�������&G��(���0�l{�]&"(�q9+t�}����@|����^a�nu4Bޗ��jw�	�����*y}e�����ӽC�H�CW���|e"�K�,ǆ�`�íN=]b~*��s�h3pX���Ь�J������pك �%�K��^/p#��I2�8��[�@���=aS�H��ݚ�Н�`&c�'N�j���$�a���NM���$f��_Ub��7��G_���;�P�t�5�׹����忔8l{�]&"(��0�"�˲yQڥ�#�Gւ�Ѓ0�ߔ�;�&���b����~�]��/�\����P �"ƾ��gx�׈�xIY��8>h�|�Ȝ��quA0�e]'\gWg��	�Z�kfc�_	�Ƽ��S�J\7lk�p�+N᢯��0�8D�r^�Hd���"sS<�0�zG�������&G��೹�C�A�IS��[;\v�a��ƍ2���l�����g�Z��3��a���!@�f")u��r��Y��8>h�|�Ȝ���q9+t�}�|#HK�� ��5%q���f�e�!\���x�sl��Va�ir&�����2q(���27:�������&2��OY�J�M����!�`�(i3�Uʮ�V(Y�t���1�g״$(�>g�fĉ>99��A0ok�����F��O�\E�W��4b�⾰��bK���żh��e� S�p���k��~��/6�o8:4�I���c�90��G��6�iI9�o«IX0F�M�sݸ�/�gxjzӝ���I(͂��-������!�����ִ���	ɩ���@|����^a�nu4Bޗ��jw�	���|#HK�� ��5%q���f�e�x��w����֯���,mk��L�������&G����l��>J��Ëf���:�I����Q؃�L�/�Ѿf��6�$VV���ݚ�Н�ٮOS���pޣHV�v&
1����nX��-/a8!�`�(i35i�a�vb�^օ?D^��՝� s�#���k$ '9�и��{.��_+��y�և@>������$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vx�6�~�q�
4������; i�V�JD�IX0F�MV�ҁGG%4vkz����`���φ��<�6�c��:� �����"sS<�0�zG�������&GU�z���K� |�>��̢k���F�KD�Vr[/}>5��0�B� �b���H�������3rnu�j�fK������&G����l��w�|l�>P"G�wk���zܳX�P��%�©p��;�{��!�`�(i3u�st����'�PD��	��x��ݚ�Н�9O�m96�o9i�!>������$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vxyk���]{�H�^A02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�D�{�ը7�<P�qb`2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �,�E�ϣ%�t�/7��[��IX0F�MV�ҁGG�.Mm-;�d=��¾ȼ\���F�`yx�>�+X�M?��y�H������N����n��>�my$�N��o�/���;WJ�Vп;3�����I����~u/��kOT=�40]���8�C�Ћu�a�E�Rq���my$�N��o�/���;#&WJ�z�6�2�^�?�/��kOT*qA����6\�4�@�� �-j�1tSjv�X19�-.|}�ڎC�?�x��w�����ԬQ����5��t��[���}��M�?L}�7�����&G�0�9&،�Zg�x��.2`�#���G1[��y�q�9�ͭ����qJt�_�/}	��n�re�.��:�4��f�i�Q2X��K���E��!��c�^[v�5Q�͍�Z%؃t����}���V|Cy�W�CbE�"��K�w(T"c!s�$f��_Ub��7��G_��:䩒=]'�Fr��j�:�����e�yrJ�āD����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc� ���j���d�a����,��y˭��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���m�(M�z}����IX0F�MV�ҁGG%4vkz���յ[+8��r$ɓǃl[�Ƶ�1tSjv��m��
��:�'�:�{_8�Y��=�}�Vݨ!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^�ґ`�g�y z�P��	���QC�íN=]b~*��s�/$�ߺ��]���޵.��6��t�b�!�`�(i3A���|��`�Y���p�_5�?*ٯ����z����,:&ȨّJ8�o�w�xˉu��r��9lD��XH�|ը�K�Q�c��~����}Dq�f�m��;���1&��*�("��X2��4�j:��e+�������� h�ҩ��m��
��:�'�:������W���b�0���Ě����E�i�m}6O�D mWN��ܐ�}�J�S�8�X ��f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���������L�Y&��m15se��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}��T1�8K��X�-�Y���U��)���Y;e�iK!���d.���8-|�D���"sS<�0�zG�������&GK��ft����Y�b�������9�ƍ2���l�����g�Z��3��a���!@�f")u��r���\!�U,ܓh�,��R��3��
�M����d��-��!g��J�s��z�
1���;#o�]�ʄǘ9��V�9�6)b!� 0/0`9N1�
�M��.��g�F��6x��w����Q�TyǨ.�2��N��-����P#+_]ݱ�m�
���nGW�:!�E�.g"UƄ3[�g�DPp��k��^�1��[��o}��MX�w����D����K�f�1tSjv�K��ft����Y�b���v�Ѭ�����R#�K�|y:�1^0lfHN��R��bP�63Z�t�5ߧE4��Fr��j#k
z��k�m�
���nx�]l�i6�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl����::R�{�>����t2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������h}�"+�{z���K�h�&~pƹR�"J�;����g��徐�ߑ�Km�?0c���<�<��(�;�n _��{�5�Y�w��i9h��W� c�.[K��m��S&ϊH��c�쭄]���Ske޸XhZ[�}Q�9�ַ���5�����,p�ն��95�2����Z�׭ �k�30: ��q�[���1x�"�Ag����<v�Y\`O.C�x��7��c�^[v�5�Z�|��w(K7͍��|��W&":�@��v{�G`,9�H�W��-���֪�K�;˞H���@���4�c[2����ZqJ*A&-�Ri�H����JAA4i1�*_k�B�a��� h�ҩ��H����ڻ�+���i��ċ�!1tSjv�!�`�(i3
/���p\"�!˥���KS����<;�$��У2=E���3	�o�{,\�0+sJ���|e"fĉ>99��A0ok�Ra])n#���r�����Jo���j� ��7P��'����u��r��!�`�(i3����Y̀�3#O�2�B���s�����X�X���`��,n��뾦�!�`�(i3��Ě�����}Dq�f���Ě�����}Dq�f�fF�5.]���E�i�m}6߸��S�Ȍ��9�ڮW;��|Bΐߧ �l�}!�#�bX�h��M���`��&0���Q��Ӏ�FQ
П�мBAϭ!�����D)���w=�ֶJ��:������TtU��
�IȤ7�����t�T�-g�
Mz���n H��èV㣅Dy�'0: ��q�;&=7�kJb�z'hۉ)��d�7�q�5�����}Y�u�U���2�B���s���EG����'g`$�Y/!���La�2U�5;����Yk��]�Q�&��H'o�a8��v��ONH!�`�(i3�\!�U��T���a��o���H�RtV�^�#�-�p�h�
d���@f5��TF ��*�S#�B+� 9>P9<���F��}Dq�f�HN��R��bP�63Z�t�	��x��ݚ�Н�X19�-.|}��FL��G��Hb� h�ҩι�+�t2�c�^[v�5�ܾ��mk�9$[{^+#y㪁��i�u״$(�>g�!�`�(i3���F��O��ݚ�Н����F��O��;b�-�2�Ct�w#��@}�	76�&�φ��<�6�aT��3G?�d���&���TtU��
g1�MVjg[:%w�&/.����#�>�n���X��RLT��T�٥��T��Z��J�~����p�q��l0����Y�)en7�F��(�[�o��_�Rv�䩲$��8��I��.��|ȃ�A(�c���_G��Hb� h�ҩ��T1�8K��}!�#�bs��>H�,b�z'hۉ)��d�7�q��k��^�1��dc�@c�����h��-�����Jo���jk���%�8�Va�ir���+1�;�.��1��!*��*8��!�qgy�`��vNd�8��k�Ss��Zf���g�F��6�	�¥�S`Q�TyǨ��&��I��"ǉ�t������z���x��y�o�!�`�(i3<���d1x��r-�T�����+v0: ��q�e>%����T+���f��,�,&��`�2,�!���������d9=���u��r��9lD��XH:�b��tv|	C���0: ��q˕��h `��;b�-�2��;�P�t�5m�ڨ�hծ��Ě���aT��3G�IX0F�M����Y�)en7�4_&��,2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�$�/T�!�'��񫯃���{S�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl�܅��6���+""�?��n��J�
����[2BĊB�#y�/&*�vW(�����bʚ���"�Ag����<v�Y\`���8-|�D b��tY������`��nF���<�W�.�P�	��
�Q�}�R'cf��!sR*��d�(���B���o��+eQL�0� [�3	�o�{�p�l�~�Q?M8�f2]�Q�&��H'o�a8�J�M����!�`�(i3i}B2>�~ �<j�"�AM?��y�!�`�(i3ʲ��U�4f�
"_��P��]�/F��?D�8��	��x��ݚ�Н� b��tY�0�����V	����/��kOTfĉ>99��A0ok��$f��_Ub��7��G_��Ct�w#��@\E�W��4b��Q+��
���t��{Ck	��+�a޵��	��!�2��\HuE�x�n���R����!k����@�=GGφ��<�6�@a� ��fFMqlg{y����i�q,?5q�D�E���'���A)�'ž1�|�'����u��r���<��a�X�r��ڵ�r)P<�ܓ�Y�̢k���F�KD�Vr[/}>5��0�B� �b���H����D3w��'��b~*��s��0M�Ŷ�Eʨ�`N/��R��3���:
1���Ư����z���܌��!���uxrBZ@2`u0�F��ay�z�v�À����@���l��[���}��M�?L}�7\���03!�`�(i3;s�e�$X�}���钝���3�#��}Dq�f�m��;���1&��*�("��X2��4�j:��e+�������� h�ҩ��m��
��>W�~����2�I�b	�fƏ���%>�rGO�D mWN��Ě���aT��3G�IX0F�M�~�eW�Ae��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!�0���ɵx�/.ؘ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc6^-Yu��_;��up�6��o�
w�f�:"�G�}��d���!i��f�,�k]�c�jd�L�\��;�,l\�=�]y��I����~u/��kOT	�%��6� ����7�*���́;��|B���o1��Ī��p1�;#��Hۭup�6��o�
w�f�Q17�b�����$1&O�|����è>�����0��� Љ��zռu��R�~�S���D�:��L)��tn�u����L�Y&~�ؤ�\��MQ���0�+ʛ�����Γ8�dKa�����Q؃�L�/�Ѿf��+�_0c ۪�-oF����7Î�I&ۛ��*ަlCi�n��Mm�:����e�5�Y�+��|T�b�z|w:R��i+��ɢm��@0�ڥ����ȾD3w��'��b~*��s��0M�Ŷ�Eʨ�`N/�xP+�L��k��������d��-��!1U��y�NӼ0��J����wg>M��b�Bϱ��>1J����C#yJ�jF�ཕu�ާ�����ݚ�Н�!�`�(i3�����z�/v7|�|��&���IX0F�MV�ҁGG`5:�����8-|�D�H����Qw�c4~Nr_�mS8<�n�ݚ�Н�	�%��6� ����7����|e"*qA����6\�4�@�� �-j�1tSjv��� л��X�j(�w�|,א�2�0��D���B�-��8�>O- GQH���U�گ x��G64����d���a�:pS� ���@h����v{:��h��x��8<�G�6�!~�#o�]�ʄ�߸��S�Ȍ:�^ao�&�U��f�!�`�(i3MQ���0�-��h��ƍ2���lĹ߆�p�h��7�^t��d��-��!g��J�s����0�|�6��t�b�!�`�(i35��
.�Ӽ0��J����wg>M��b�Bϱ��>1J����C#yJ�jF�ཕu�Xt"�K�AԢ�a\�'QZ˂�b�Z��M��4k���r0��K�Ǔ�\� h�ҩ�7�wtMM��6�a��״$(�>g�
�:qEp�;�P�t�5fĉ>99��A0ok�׹���C���N��zL����ڻC�i�;��|B�:�(��?#�ˏkY�J+�WTIM�,!hޖ�A$�P������5d��n4s1�U��B��-_S���\���T���I9���"sS<�0�zG�������&G7�wtMM�P��ì/��kOT*qA����6\�4�@�� �-j�1tSjv��x��8<�`u0�F��a�Va�ir���+1�;�.��1��!*��*8��!�qgy�`��vN1tSjv�7�wtMM�P��ì���NM���$f��_Ub�F�S�1 ���V�v���4N�J�ף������&G��+�t2�T�3�7�*l)P<�ܓ�Yfĉ>99��A0ok�����F��O�\E�W��4b����A������f�6�H�^A02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc0l)�┗u����p����t�T��?E-h��`f���sd�G}%����3fX�?���'�V�2�~ڦ'ž1�|�'����u��r����~Щ�n��뾦��߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#���N4�>y�pA��M?��y�!�`�(i3�	�%1A��b+}y[HN��R��bP�63Z�t�5ߧE4��Fr��j�p���"[(�i�x�n��{"[)�`����ǆ�S���Q=-C ��U�