��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��]	h8��`��(	�t�&�u�"��U���T��ײ2��>���^k�/7�?1�(�c��ly[�$D֍C95^T��#� _�_Ü�@�hF��W��`��q�©��ല���?�;��XC:Ҹ������b1Ø^���#K���lӧIA�a�V��R�}9����D~;yJ�'�دv)h�V~�$v�p��"}�v\-8�������>�`)���a��rl�ʩ{�Bf��� ��|4�VDG+�������X".��>��'��E����F�Rm�I�|^�Q�;(1Z �bRw�����IL�+�{Dr[��	�� '�T����g?�J����m�Q� C�-B��<���2O��'HY-��Yk"1/�p�r�ɹ���� �]��;�I�Qg�@zh�S҆�|n����Շ_ Q �y�N��Q(�V͆J�Й�m��x����y7���̖�}�Ϫ�h�C �@nk����k�&�J���qݣ��6Q�eѢ��x��!�v�j�|�㈱�U^��\�4�s��{��]Qǯ������W)����VIW	I��?G�~�MUs +������\���T��U	�1�_u���*����	�����	����LO9� �Ŭ��2Dm�x]��.] �'9�����L.��6�H�.���2/�f��=V"N�^{")8�*I�ց��6 �����Y<�zd諒~����L.��6+Q)?^R7D�y�B.h�hC���(:�J�5`xt��R�/E�CԵ�_�!���<< �sN۪�c�	u�~Rp�,k���%k�&ָ��sE��D�őⴔIꈸV�MT7xB2I�d�HnULkIh��:h
�[ϸ��W�A��S;CM���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc(#`��Gcp��}K��f<�,=K�F~�?|�[_X��ˆk�=�r���x�i��p�7��Xi9�
�ѹaB��Q�//?�s�m/C�N{a�9O!JoE'U�Y�y��
r�)�Y¹w����i��T!ix�AH�k[�^��_�0w�T^�W�����%3?���kW���;��sD���L�S5H�j.F�QSjl�g�L�Xڈ*-}|��ι%9��oGo�Z�J��ݪ�nP;���7	�\�Z�م~09h�i�k1i�f1?�6K.�ُQ�����0�ea�8���`8��xS�^�����������,\ަ�It�k\,آ(&l������ nU�IÙ=�HF���m¡p~z�r,i��i���'n�^0o<H�-��*����Kp&�@���k��JHn��z�_c)���8�+�p}>&�&i�A ��E+���XP��Ȩ�wl��h�d�uY�ة�ʐx�?�'n�^0o4M,������2��̪
)\Y��7�ܥ��2��
[���p? E%n�/���i� � �	{����0�&�ͭ!�`�(i3N�By3��<�]�!����M[��Ǣk/�z�xEQ!�`�(i3c��Et��q���U�&��GE<�!�`�(i3Y%T��BPe.��xu	�>��l%i�-��TBd��pS�*;q܄}͟PP��Z鎬����
C��8q��f�kN�ı&l������\�*P�I7��-5��6��	���`y���db�\EX@�/�M^��Hm��e.��xu	�n�-�6��
�jW��D���M��ҹf�f3'"�C�ף�;�¬pX��g��U-�e�,���6+�+�uB;y�L�6yd(��(�
t��Y�{'%s�[�&B�踫g(�r� k�|6�8j��RO�I�1�Z���=�"j���b7xY�J��ev�mS��0�-����#u��Yk"1/�p�r�ɹ���� Wa�b����y�E�nwE��S��}|��XH�����,>$+W��� j�(����5�:n�|����Z=%�	���,�V`�Pt�e'J��x'[{����n�4�c_����+#��.X���*"v%)��Qcm h�]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e���b P]��i�"ٷ��	N^�U��J��"ї>п�p=	�˳͠m�xW��9u$d9�cx�S�����S8����ٺ?�R�^Ƒ����"X��[��Q[R�7����$�1i���"<璋���n�4�c_����+#��.X���*"v%)��Qcm h�]�!��	Ǹ�y85�b�
RaiK�;�¬pX��g��U-�e���b P�։-�.l?���oD�fmc^���Ф>п�p=	�˳͠m�xW��9u$d9�w�"�HߢI|{�0Lʡ;�¬pX��g��U-�ez�r�6��DP֞ �����Ə/(6>������rix'f]Q�I����踫g(�r� k�|6�8-+��B�Gݓ��E� 7�J�[�}��s�e�2l��4��a��se�ξ������ei4����/����DP֞ �����K4K�)s"���݇�T%{�;����f�kN�ı&l����[}�@��L�@����gG<D�n:3MS�*;q�/(6>������rix'f]Q�I����踫g(�r� k�|6�8-+��B�Gݓ��E� 7�J�[�cd�b����H@H�֦g�㎏qló��@d���/��=��K�R�hE!3�͸@����gG�r�I��!�`�(i34K�)s"���oD�f%g4���r�<Uee�,�Aٺ�H֞��Tj%�A��N�?G%Ǐ��� gWVbT+zv�؊)�x��$1&O��P�/GGb�|2;$�JأͽgF"?��иܖ��%����8�?�d���&�{��؉j�����t�T��?E-h��$^(?��"��h��w��յ[+8����"sS<�0�zG�������&G�wӨj]h��_--���g|�m�ߕ�E�g�������(ӈ���m�r����ЈH����@�/�M�k��G<Y�dN�<@Iv��nt=:��:5A��pt�td���5�k��^�1Aj��t�35L��$
8��2�ֈe�cN�0��ž�Ć�T���7X���c�}��
�t��T&���LQ�/81tSjv��wӨj]h��_--���g|�m�ߕ�v{��lw	�����4�:5A��pЈH����@�/�M�k��G<Y��������&�G}��ݚ�Н����F��O��;b�-�2��;�P�t�5W?�;�끣�os�鮊Vo����6j�"Hs;&�C�����#;�A��A���`����oȺf�畮�e��d[?�d���&��ꢤ�Og>ݣK�6<o�����w�_--���ggO��;�3t 7�J�[���R��u��g��L�,�ꊃ_V��	��y&Qe�}�!����ݐ|
���혅vº�w�⽒��8�>r&�,�Aٺ�H�f>x�:	�W+��W��]G�ߕ6�o8:4�I���c�90�Ǘa��xO.C��|#HK��A(�c���_G��Hb� h�ҩΤ/�cLb�����صW�my$�N��o�/���;�Ra])n#�璓�c�������t �[l;[�G���KlG%��`��ǚ��ظ
��@�U#;�jmT�#�,l����M?��y����Fz�΋O�»%���]c���HE4SG���Z����Sz�����!�`�(i37�A��\R&k@C�Ɨ0z�cUL?��[[�L�1p/-�������?�/5��"}�a�x�mj�B��Vh�EtC�<��R@��"�!�`�(i3e����R,�!�`�(i3FwZNE�&tS�D�'���Xw�j�7��AԢ�a\�Y��Pv����ʗ�%E+�}��D����0�� 7�J�[|�m�ߕ��[���#�!�`�(i3�5ߧE4��!�`�(i3��4-�c�{I��L�1p/-�������?�/5��"}�a�x�mj�B��Vh�EtC�<���v�9��HN��R��bP�63Z�t��Ě����E�i�m}6߸��S�ȌX�f�βB�.�g3Z�j5�{�S�g�E8�W�~����oȺf��A?�87U�?�d���&�_|�9�0ݤ|2;$�JأͽgF"?��иܖ��%����8�?�d���&��8�c-~���bY�}��φ��<�6�@a� ���N���Q'݀�=�յ[+8��H����Qw�c4~Nr_�mS8<�n�ݚ�Н�{k�h�+�=<�6>e��0�U+�qbp@�!�`�(i3�Ro�G/]%�z�-uͺ�s�η3G��Hb+�����;y��v��\���
^�ݚ�Н��
�t��T&���LQ�/81tSjv�!�`�(i3DN��5\���51�X�c�rs�i��L�������y��!�`�(i3��Ě�����}Dq�f���Ě�����}Dq�f���ܐ�}Ęs�WGqD7J��0Uw�R���y@�67d�aT��3G?�d���&�	0vn},5���}�$Ɍ�D�ݓ#_}p~z�r,[�?��{W��d���!i�P=��1�(��`��&�u�Y�KG�	�v�3� k�|6�8��:�EB�Z5�O�%E#Pq�\E��0Z'pǘ���Z鎬�������(���fD=����e$r�t�}iV��	��yO��aQ'��^�%�P�m�V��	��y�q���bc�ya����6�6����D5�|أͽgF"?�Q��ǺΕ�f�f3'_��s�֙R���Bk�d���H��H�2��z�b�4��Ǳ߁R�^Ƒ�өwo��Z��Ac<�p{�5�O�%E#Pq�\E��0����E�I~�*0�ŷc?KYC'v�����G eK�lݧ}�	76�&�;��|B4<d��
~�_��.��ϕ��q�"��Jl��q<uiF=�xo�R�^Ƒ�өwo��Z��Ac<�p{�5�O�%E#P�G�dE�h����E�IȪG:vmX��u��g��L�������<�^._�}�	76�&�;��|B4<d��
~�~���.�;��|B31F��~Gf��x��9�Mgw�� 
~�F�,���XF:��GZ>.�0����ڀS��d���!i��x��=;Y�ۺ�Ub�!�V��u��d�uY��s�N
�u�}�T�\ ��;��|B���r����+�uB;y�XNAA���v{��lw	+z��D�H�}�	76�&�;��|B�T'[/Ʊ�&UX�{6j�"Hs|��^�p!"���(�e�Aa�R�