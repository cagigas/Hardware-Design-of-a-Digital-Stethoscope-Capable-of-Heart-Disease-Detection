��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��k�	G���%��%���UQ���?6U���T��ײ2��>���^k�/7�?1�(�c��ly[�$D֍r�	�tX�)�`���$��[dm��+@ˏ^ow�Vx���_>{������6��H4ٳ�k.w�.u���ŏ|{T%�at�3������ͧ��G�]�ڶ�Us�JG�DGsc2�aB�>�;�C�l�����h?M����bÛ�>/�F�q�\�0k�5k��J�|(���u����l�|���j�I�?g�f	T��i����Zߧl4���0�?�1~�x�cX`X�B%�r���7�8�.��9����/�k���hoP뫼b#Ӡe��?�F��&4%�}|x�el���7`ɝ��kN���9�ĒTC��0��`�R&.1�w��-�95�]����k?�w�>��S�@~�w��!s.��"����dLC��%��w��^m�!=�y����h�}T��nJ8�8Y�&�\�#�W��a��#�Ԗ̋�N�u���u��Uy�PD4KU7B�����<�[0YY���\�4�s���rH
>8Y�&�\�@N��B@B����n;�q�m���mi=��B�-x=�WD���4B'���S�K��i|ٓ������v9{�$W
?%x�+�� fג�� y�dH�]��/�2�-�]?�B�nI�4q�Qt!��c��<%>ì�oJ5�%,�k�W��T�٥��T�Sҥ��|E�EYZ/� c��(�U����	x]�����O���8�t��s*ո{�x�G�F�����OwꅂF�-!d6߿��b��'�� |X��M��"�D�u���lٽ�G��k�8���҆�|n���u� �(���jV%[&��\�۱��ѕ���Z�[�0�7٢z|Mߘ����g�/@�G��P�?^
ر��ZXty���`�c�~e�0�We���ܮ�c:��1��q������-i����^!`w�� ��A�]�B=>_�o&�8��/M4#>Y��<<�٤:�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��r�����A�F�7���3�GXS����E@��~���($�J.���
�=W�֯��i@F�5�=h�GD�#�̔"v��ƒ)?˳R����.��ѬL�1m��+Y#_WӢۉ���2=�l�����뙇�� E���Ӿ���	���qk�ZV"���:��#tCE8�^��������3�C�p侢����U���h����S��i�twJ:�FT�c�$��b9���1��]2�?V�Ľ��'�\�nﮅ���gzL͊�q���1m��d+0�l�R<�q��f�}��h�'f R�E����F��j��\w��0]��0�&�ͭ!�`�(i3c��Et��q���U��>�w�Y�#���@d�E���-��%M�rs�i���`�M�	=̞��>����� +'������݃�Q[R�7E[��\ ��;Ai�Ő��-��%Mό���.Ӂ��̰�!�Xy|�W�����
L'���Xw-�}��dB<�L�V_N�By3��<�]�!��	Ǹ�y85��ٍ��%ڞN�gl��ܬa(􆿳����^���(R\֎u���sRt�7G#+��\w��0](@X~�H:�W��7=c��Et��q���U�[��N���v�Z�]2�y�Z鎬�����	�7 �#�\1^O��0ˋ��I��w��,>����C��(R\֎u��ԟ'�D�7G#+�Ǘ0z�cULjaGkƊ~8����\.W^�V]��}<|������N�?�_uM��y��I�+��T���jB�Fg�Y씤`��p}RQaI+اy�TՄl&K[�
C����[5`� Oag�qod�֓��+��T���jB�Fg�Y씤`��p}RQaI+اy�TՄl&K[�
C�m��P��I��'����cԱn��aМ��IÙ=�H�R����/�R�|_v�:��j��ji���+�z�m_ �e�12R��Ûf�̅J�9h��$`3d�>?�^���_�b!��u�D��ɍ�٠�и�0�G�w�^>��p3�+��m\���_j���5z����k;{�R5�5����n9�u�#�$IX��V̇���˳͠m�xW��-#��k��b�`3E��Ҷ����2E�$��n��:�n��,Nzm)�W+`�x�o/��A����~��yZ鎬�������(���pl!�6���;b��g��U-�e5/�=��kb!��uፏ����V?ː���T[���h^�+�>8
�O�t���o����;�Ӏ��nrm؊(��@����gG=%� g�Vv�5)��Z^7s�9���o>��l%i�-5�e`��9�iK�D�b=	�P�g�Z鎬����V��J��3qE��6I&���#��1 bL�o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc?��΃����7��Q*p_�ɬz!�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��OC�0M�|a)� ����35}jds�c�w�",oMG~�K�3�Ƅ�u",oMG~�pm�#�ŀ��v;N��-2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR����#�ͩ�n?g���3������$�c/�M��lj�K��5�ʏ�F���ٷ#J�C%o��T�
g������:[d�dݵ���n�`������s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hMQ���0M�,!hޖ�A$�P������5d��n4s1�U��B��-_S���\���"2�HJ}�r$ɓǃl[�Ƶ�xm��s��ݑ���&�d�����lɢm��@0�ƍ2���l�����g�Z��3��a���!@�f")�j�&�-*�c5ew�|�;�Ojz�$�AՁ�Va�iryP��C��?�T'���̻���S��!�`�(i3fD��j���eK�	�$V�#o�]�ʄ�;4�zu%��XW�G�<b~*��s�
�I�b�_F�1tSjv�ݑ���&�d�����lɢm��@0��?D�8���������+�t2��iK�D�b=C��CFv$���b+}y[HN��R��bP�63Z�t�5ߧE4��Fr��j�p���"���,�֎�B0��5��Xy|�WS1�ӿ�Q�ЙMǿI?��m݊#V�Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hKp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>ha=�T;��W�.��A$�P������5d�	�+�&I(&�L��'ž1�|�'����u��r��'V`��bޞ�>��[V����@|����^a�nu4Bޗ��jw�	��x��7��74/�����w�`L��t���Q�5ߧE4��Fr��jL��[��M��qx ����	+��g��=R�������泞Wacʞ�Ck��N�DNlF�{T�ō�恇wv����èV5�v��cg7Ԝ7(u�/�"����N�PBaE&U�)j�S���ܚ��@��f�\%����e��!�`�(i3��_	��Eʨ�`N/������&G!�`�(i3����-J2�բU�?�2h��艅�%>�rG�@�	����ʁ���MյFr�S��PL�3��Y$�VZ�ڋ���Y�ُC�YH�!�`�(i3��_	��Eʨ�`N/������&G!�`�(i3��B/�)����bX�'����u��r��!�`�(i3��w�`L�U5���M���[ӝ��o7
�:qEp'{w#/ B!�`�(i3��w�`L�U5���M�����yV�a{
�:qEp�;�P�t�5
�:qEp��h�8� ��0�|��';��#j�ݚ�Н�i|�rBY���N�DNlvr5�Dѯ���-����!�`�(i3�FW�DVx>74/���1�L�3�!�`�(i3�5ߧE4��!�`�(i3�5ߧE4��!�`�(i3/�"����rE�s�Bv�K��ٳ�jCH�d*��=����h�qB��S)��}Dq�f��\!�U��0�|�_�mS8<�n�ݚ�Н�i|�rBY���N�DNlvr5�Dѯ���-����!�`�(i3�FW�DVx>74/�����ǔ�-!�`�(i3��jVѭ@!�`�(i3�FW�DVx>74/�����`V�6�!�`�(i3���F��O��ݚ�Н���?2�}X9��|��ֲ������ h�ҩ��H����yP��C��?�T'����������ݚ�Н�jCH�d*��=����h�(-���[���}Dq�f�՝� s�#���k$ !�`�(i3����-J2�բU�?j���4(!�`�(i3�5ߧE4��!�`�(i3�5ߧE4��!�`�(i3/�"����rE�s�Bv�7: �"~*jCH�d*��=����h�'i`.���}Dq�f��\!�U��0�|�_�mS8<�n�ݚ�Н�u�RV��,��-G̙� F���ضo{�U���<�����Mʠ�@I���w��[#M�=~~*5�tD�#k0�!�`�(i3���L2��AݡٍTZמFS���E[��t�9��|���5��<�>P�"ѹm,�3�(J(��fh����爮��J���ݚ�Н���?2�}X9��|��ֲ������ h�ҩ��H����yP��C��?�T'����������ݚ�Н�jCH�d*��=����h�qB��S)��}Dq�f�՝� s�#���k$ !�`�(i3����-J2�բU�?���~t�!�`�(i3�5ߧE4��!�`�(i3�5ߧE4��!�`�(i3/�"����V(pyL0DMlE'�! CH$�I��*�M/*�3҃�q�}���}Dq�f�ppE�"f�Q������\E�W��4b-Ukc��Rg�a%�}�&E�*f*�(4	d��R�w(�|��`p�~(�M��1�, �F�̃��HФ\�g{I�"�on�~��2�>޶�[��o}2?�;Ȟ��
�Iӆ��c����jVѭ@!�`�(i3!�`�(i3v4{��Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�(}�����#`7}"�}��O�l�<P�X�۹hDl���YKp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�9����(M�,!hޖ�A$�P������5d��n4s1�U��B��-4��)'�����u��0C�r$ɓǃl[�Ƶ�xm��s��'9�и��{4hz�<Ρa�E�Rq���my$�N��{_8�Y��=�}�Vݨ$r�t�}ik+Q�h'�Ȝx�5W ��̫(�H��
J��7�:t�?S/��ۀN���o�u�/ q��j�J^���c!�}q���f�e�x��w�����$J�L߉����n��<f���=m�n�V�EVt�`t!�`�(i3�!���MEʨ�`N/�<<��lp��N�DNlvr5�Dѯ���,:&�fh��[�? �e6j��9��ݚ�Н�7��u������v������f!���®�b՝� s�#mݹC�ҩ)����bX�d��-��!�$g�ޖ4���(;���-����!�`�(i3�����V?�k� ��"�?��۳lU����Ga�Jv�w˅(oHN��R��bP�63Z�t�2�2���'���r���b�����¡����"X19�-.|}�íN=]b~*��s��(R\֎u��Gj7�uz�gVdxQ,��[��o} ��:^"�x� h�ҩ�'9�и��{4hz�<Ρ�cl�j�pॻ}����}Dq�f����F��O�}�	76�&�� Ӗ�t$�)�vxݳcF����0�"�˲'�ZX^�O�<�Hԯ�!{1�~���W�3�-8y~��׺�o��_�Rv�䩲$��8��I�:Fa�7���^�#�nish�Ž��2G�,��R(bs��2[�a��o�����]�KS�%t̓�@���'|F�{_8�Y��=�}�Vݨ!��"� +}0�ʂ�j�Ï��	�l�lM�3 ԫ[=�.n��:咦9��0�|섃Va�ir��[��o}�+��8�T�d��Ɩ/ ��Aݡ��d��-��!��KVט$�W��7=#o�]�ʄǬ�$gQy�f�ҫ
OԐ��-������l�^!�%��ږ���⣮`��+�T[n�߆�p�hؤ	ͰZ����XW�G�<b~*��s��[�#�����?ln`E�p������(;��B� �b�й�+�t2��#✲�@��kb- m޺�����9�<F3�@�@W���%>�rGO�D mWN��Ě���aT��3G�IX0F�M%w�*�7��q�3� U�%t̓�@���O|���p�@OM.Ir{U����ƽ[Gʜ5�1���~!�`�(i3��7I���Y;�e�O�!�}�Ͷ�,*^���H> �}��%v�\����U�._�AԢ�a\��$p��̧+ڰb��Ƽ��r����!�`�(i3v4{��Q� �_ttbh�m��d0φ��<�6�@a� ���N��ȥ�n4s1��7�癆cgQw�c4~Nr_�mS8<�nt�{#	�x�u�#�$IX�]�p� ��߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#�(R\֎u�eK�	�$V�#o�]�ʄ�;4�zu%��XW�G�<a��o���H�RtV�^�_��*��j ��b;�(���27:֭��� �*P�엫�u��r���2��}���'��L��K� |�>�
�:qEp'{w#/ B�2��}���'��L��v{��lw	���l�K�F���m¡HN��R��bP�63Z�t��Ě����E�i�m}6�@�	���Ĕ׹�S�C��-<o�;)�yԸڇ���<w�T� �f&���#��D<V�-�b�+�