��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�>���U�_�4�0S�����xnP;���77\F���r����&$9g8�M>PFWD#�z":���ӳ��_}��0w�\1����K~�j�k��� �Pq���Ɽ�Yk"1/s�\"�����p"�+ڍ�P��*r���`���N�w	*D���y&�f��+K��[y��ڂ�Vs>�+���,>z���/lt�3� P�;��1�-��⫯g*P(�C#<�:z����uP!ߌ��˼�{�&���7�os!w����]��4�:j�l�,9����=-��Ǘ��p��W*[��HMiL���om�Q*���T�K�MV}xj\�iW�(� 0�D�A~����p��ؚ�fD�~����pn��-�4ڭ	���
��M!�nz��m��+���J q�v����6��w�1&�u�"��U���T�����\�4�sW c`k���(�Y���mM+­�\��S�Q�L�����Y�b�Cj�,\ަ�It��vȯq�
� �AH���g���	�'�Wا[b��(�s�J�=�ʝF@�4%���IR.ux'V�vЊ�[-d�x�����q�M�40�W�wƼ�{�4��W��#0��<JTT*��@n���SۣFߞ��G�٘�`�Ocᑕ:�,��JCq��jr#�9l$!kdq��]x��	�VE��t����G�٘�(�����3Y&{ �ŠB�N�M2rӪ���!�Aͧ�	&�~��FjrHS�w�MH��j���r���+W��YJt�,�y"r� J&g~���c*& z�s�ђ�B�~f��0(�/��$ }2����T���Q���!i��ӯ�02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vce��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�׍E�+��
���*,f$�7Q0- ��Ck�fÜ�2/���}����сsU%���n��/���Û�E�tw:g?�y��h�I����uk1i�f1?���b1�F��,��n�2��C�`Q���Ӿ���	���q��q�©�����<�������~s���^��	���,�V`t�iZ]XF��������;-;*�7����]n��,ԯ���gn����fԱ@j޽���Ǜ�����������i�jݭ�F����QI�D/����ʊv.s/�B{�o
��ʺ�;[��#�ڊ<?@��[	J��;ι��QG�����U��!�`�(i3x�]�V��;���Ӧ��S1�����)��j)yc�n�.�_�t�7�ܥ��2�΂��F�V��Q�S���>$T 
����>s��Y�&�E����F���8�TP��������ERF�G{؍��R��j�.(Wx*9��?xs�S��'�?�]�!��	Ǹ�y85��1}�\���;�¬pX��g��U-�e�,���6+�^�9.�JQ��{l�f|��rs�i�� ��*b��0��E|�,�CyW�f�tR�wX�Ռꢤ�OgI`H�S���]���c�A�L'��!�a��5�%]���a(􆿳����^���`��׊���TD���rs�i�jf� l�Ǜ������CyW�f�tR�wX����d\��N�By3��<Z鎬���������o�	����}��S�)37J*u>����CΫa������<��z��}���w�V�"-4��h�]8+��T����oGo�Z�������/�)��ɖa�\7�"
qWa�b����y�E�nwE��S��}|��XH�����,>$+W��� j�(����5���ռ�j����)w�n��ukh���9tf<[f�c\?k%���ۂ�3U�?��)�Rݛ��%�5��lW0۳�*ȑs;��|B�R�.6�W;��|BK�B�<�t��I%U��_bM+���C����
&h���ٙ���O�Q���*��P�Vr���F�!��c���Y�҈�FQ��ݢt\�y~?��t�iZ]XF�hx��G��!�`�(i3�v1a{J�^�|n�M�!�`�(i3!�`�(i3J�]�RU�`���!�`�(i3��<E�f�y�-
9dZ��|�H.z!�`�(i3�;�����^��&X!=!�`�(i3��<E�f�y�-
9dZ�
I�Vd��!�`�(i3�;�����^��&X!=!�`�(i3��<E�f��V�mK�b\��Mh�!�`�(i3�;�����^��&X!=!�`�(i3��<E�f��V�mK�b6�X�$�!�`�(i3�;�����^��&X!=!�`�(i3��R~�e��ד*�h��F�v�C!�`�(i3�������a�_���!�`�(i3�Z�r6�ԙ{<qH�~�!�`�(i3!�`�(i3J�]�RU�`���!�`�(i3?�ᒹ�G�!�`�(i3!�`�(i3!�`�(i3rQ�4��+��S��?�F�`���+�r'Z1p8��e�j�!�`�(i3!�`�(i3�&8�,���	ǗP؊�á�~O��&�C�/�<�W������!�`�(i3!�`�(i3-��U��p�K�{R�^Ƒ��f�?ǉ�="D�
�	+/O�Q� !�`�(i3!�`�(i3�X;p`�Pm~�@P&�#�|M�d�>b�eIG��Q�q>x�-#F\eڲ!�`�(i3!�`�(i3��g��E��� ������$Y� 2��4����7
!�`�(i3!�`�(i3�b[�u2�G�=����ڄ������b�Xϋ?@,�Xʚ@h!�`�(i3!�`�(i3fC��T����ܼ��]"danS����˥����AB9���w�!�`�(i3�#�q<��8���_�[�wbk�$+��m�yo���|��Mb��y9xO�`G��
��E�^��֯b�jT�.���ܴ���~�Y���(�}�Π�cC!�`�(i3!�`�(i3!�`�(i3B�O�%J(�
�cc�V��ݚ�Н�����o��,�Xʚ@h!�`�(i3!�`�(i3�AQ�0G�F�r�f�t��5Z��~�Y���(���;����f!�`�(i3!�`�(i3!�`�(i3�F�7��Y�
�cc�V��ݚ�Н��#�@�o0!�`�(i3!�`�(i3!�`�(i3X&|a�#�I7��-5��5Z��~�Y���(���8���g^��/�d!�`�(i3!�`�(i3lj�w�/�e S]#�e����kn4@Q�/�!�`�(i3n&����_�a�/!O�f�?ǉ�=���&Z>0���oC���\�tP�;�s�٩��� Ī��(�����SƏw0�����
{��{Z�{0�;?\�tP�;�6�5�p���g�+��.��	�si7��ݚ�Н���O�q�̍�����Jw����fG�E
b�+|�&8�,�oٸ���!�`�(i3��/z*x�n;��|B��)���i��q�#��3Ah	)ޟ!N�'�y�G