��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��maC�S�s�KT�=�]��;�Iώx�t���E�L#uc��WŬ�+�-ޗ(huUPc�k�u�}�FNy�N�H�d�j�m��+�Ƽ(��hl&K[�
CN<��;��� B]�pE���	x]̃Dj#^Da����M�r���
�'�ө-$J�z����)�,�˛D��w���旴4�����:��@���b���$[+r�bH7�D�C|N��^ �}w�*.��>��'��E����FDR��f��Us�'U�?K4��G%�L���om�Q*���T�K/ZT�@�t���@H���n�GE!���I0�������p����̴jz�ҲȮ$��fb���z�������@����9^�"nq���z!$��R�ǌ�꟪���K� w�;�d���N�tכ݁=9�|Z���ߐ'�[�Z���1VU���+L��h��X�vB#|y{����P7�.yt�gU*Z9B[�^������+�ͫUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcMD��y�sY2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�#CC1X�G�ۄ��O���azhݪm����Y�{'%s#K�v]|nf<�,=K�F��N��j��D���s���ئS��.V&��B֥��f���F*�#C(�����s����Ct�z&��ÃlO ܅dxF���u$J��<
DN�%Ah�%4
>��XP���C�&NJ=رx���9pk�o��jV�{+��]n���b9����$�n������ л�A�.�hQ3'c���������n|���띂ii�4];ˍH����Ү���/^�yQA��c?A���$v^�1�N�Ae�#�k/�z�xEQc��Et��q���U�ЂDa��(;�A)k�e.��xu	�>��l%i�-��9��稕v�ј�"��Z鎬����$oi�~ƴ<�6�Q=j���$5�?� �٠Fd���e�ш�_(x��`��|g�Y�'���Xw�j�7���(}y���CyW�f�tR�wX��q�\E��0bq�Z��T�I��w��,c�A�L'z��0N�7;�¬pX��g��U-�eE������(fx��V$�w�I�?g�fl�NAS*����*�H�an�]��z= Oag���:tӫ�C+��T����~��@�.��#=by�뵵�
{y����x��F�U| c�]h�G2[�4��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��!$��R��zC{�N�ٜ2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ��؜�ۇ�|�uD��πx���"x����O�g)�X�cb�M���Z��d�G}%��Ď��J�Hmiԝuڎ�W�ҩE�t
]��v�7]�W^@��IX0F�MV�ҁGG�.Mm-;�C>��Ӛ��S�J\7J{�#�R ��Ƿ��;���Yk���'ž1�|�'����z.��W��!�`�(i3����j��3���B[=����e���A��s�R�b>3��g!�`�(i3@ E���߂�nF���<�W�.�P�	��
�Q�}�k��^�1��dc�@c�����h�'�ɳ��<�6�Q=��ž�Ć�T���7X���c�}��
�t��T&��ۥ`�M?��y�!�`�(i3D�wP�/�w��i�Wg�<πV��;�¬pX��g��U-�e�(}y��YmҐ��*V�M��nD�ݚ�Н����F��O��;b�-�2��;�P�t�5W?�;�끤g��ޏ�LԐ���D��L���p6j�"Hs~1>��]��(����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}ږ17��_>�w�hշ���+;J�@�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcN�H
��e�9X�a�}�&���m��y��(<�d������\�*�c��S��7ܪu5�O�%E#P{y����M�V<�'~1>�����#�$'7�T�f�Ǌe|&L� �IX0F�MV�ҁGG�.Mm-;�C>��Ӛ��S�J\7J{�#�RR���;h�O�M���K�r$ɓǃl[�Ƶ��I�q����!�`�(i3�� л�4�>������9�@f���ʦ�/\<���tݻ�ݚ�Н�p�n��E�g�������(ӈ���m�r����̢k���F�KD�Vr[/}>5��0�7<(�lb����y��lD�7m�T��Ʈ+ˀa��z��2�,�s�Yls�<Ԍj��_�mS8<�n�ݚ�Н�{k�h�+�c����B�:ychR�^Ƒ����"X��[��!&��F����aR�!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��jJ{�#�RR���;h�O��L���p6j�"Hs~1>��<�땮�8yKp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h����	v��(�AXP�7�Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h/�۲����mqf�����n|�p[Y���"���E��g�Ӣ�:�n*5�����e�`���;��|Bd~TK�c�i��3��^�U��)���Y;e�iKI/B޾PԐ#��go`iI9�o«IX0F�M)�|���\���F�`yx�>�+X�[�G���K!�`�(i3<�6�Q=��S<����K��!L��3w #�T�Z��&�2����D�wP�/�w{E��7ue��0�U+�qbp@�՝� s�#0�ʂ�j�Ï��	�l�lM�3 zM#��m�.�
9� ���(ٗ.;���JTv���H����o�γ�ha��o���zM#��m�t�td���5;�jmT�#�a�x�l?ud(�F�\P��51�Z���=��|+S�myu��r��!�`�(i3@ E����̷_��yC��S8�>c��6/{v=~P0:Q+�3yK������v�h!M�T�ĥ��P�7� �:5A��p�Ra])n#�vW�|�Z�d-�~E�[����b�U6�bL�s�N
�u�}1tSjv�!�`�(i3p�n��&k@C�Ɨ0z�cULE��K3�jާS��m��X�����j�5�%]���=���B�u���P�7� �:5A��p�Ra])n#���r�����2��}��e�g��)$��K���fU����z~��6��	���`y����ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6�d����%�х.�g3ZrZ�0m�\��f�P�V�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ�/��KJy�Г*9۽���cX��⤹o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vct;��C��� �R��l�&���m��y��(<�V�^�$��.��ϵ-�`İ�7�#�@*5�����e�`���;��|B�g�l$x�=ys<�+B�v��[�V}�IX0F�MV�ҁGG�.Mm-;�C>��Ӛ��S�J\7fF��v��FV��E�9�H����Qw�c4~Nr_�mS8<�n!�`�(i3���y��lD�	Sz��
�GBQQY����#H�Yg�yi��v��BPlLO+{k�h�+xއ5����K7͍��|��W&":�;b�-�2�k+Q�h'�Ȝx�5W ��̫(�8�u?��IlG%��`��ǚ��ظ
��@�U#;�jmT�#��"����G��Hb�8�u?��It�td���5;�jmT�#�a�x�l?ud(�F�\P��51�Z���=��|+S�myu��r��!�`�(i3@ E����̷_��yC��S8�>c��6/{v=~P0:Q+�3yK������v�h!M�T�ĥ��P�7� �:5A��p�Ra])n#�vW�|�Z�d-�~E�[����b�U6�bL��R���~���-/a8!�`�(i3{k�h�+,�NQ��.Y�{'%sk����w�;{�'8{1�']�JN�Zm1�Z���=�K��0Iw�U����z~)���	6�!�`�(i3��jVѭ@!�`�(i3D�wP�/�w��i�Wgd��⡙�5�%]���a(􆿳����^��
�:qEp�;�P�t�5
�:qEp�;�P�t�5fĉ>99��A0ok�׹��K{%�Y��y;�`w�R���yB9��:܆�eגb������s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}ڲ���]�&�� ���|�nKB����	�է��K�J8���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�y
�C��������,�+Ώ1;��5�}�]���LVm����1��ȵ�K���'b!��u��	O!S�E�q���U�!�`�(i3���y��lD2�û����b�N���޾��(����T�G���T׬xay�����+�^��BY�B�3�&A��S��~�r��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ƹ9��Pd�B�\��� T�j˩���	�������s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�
A�"j�F�=��Y�$��L%�G�b�gL���l�5�%]�����2���DB�*{����M���o��_�Rv�䩲$���dS@Ɵ�od�G}%����3f��,�ib�2���Z�[�[xjzӝ���I(͂�'�ɳ��!�`�(i3����j��3���B[=����e���A��s�R�b>3��g!�`�(i3@ E����x����E2b�z'hۉ)��d�7�qĹ߆�p�h��d��JXl'�T��~��?u��C@<�6�Q=��ž�Ć�T���7X���c�}��
�t��T&��ۥ`�[�G���K!�`�(i3�k��M�=q��m�3<��~�
]^1tSjv�!�`�(i3p�n��&k@C�Ɨ0z�cUL?��[[�L�1p/-�����:�(���lC��U>���Y�zb����ϏQ��8'嬘�X�h�����,H/��՝� s�#���k$ �wӨj]h�7M	�\�=��Y�$��L%�G�b��6��	㎾��;|�5�%]���U����z~���D)9W !�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��j���p�@ �P���l�0w�R���yh��7�S+����!;%2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ����#}�Σ�è��rTW��@!�|w�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc;�v�-:��%.�`�o���8�8e[m���� K���Z/N��v�qL�4@t�ޮ��ǋ�n`5�fK�3L��'9!�`�(i3�� л�iS@����n4s1�+��uK[Fh��7�S+��1ӆ�@���l�����G���5�%]����Æd�Mw[�f?�M�,!hޖ�A$�P������5d�`UNP�N}�m��{���q0�/)ONcx�:2QYeƈ)P<�ܓ�YO.C�U��B��-{��N�iI=\M��G�\���F�`yx�>�+X�[�G���K!�`�(i3<�6�Q=��S<����K��!L��3w #�T�Z��&�2����D�wP�/�w{E��7ue��0�U+�qbp@�՝� s�#0�ʂ�j�Ï��	�l�lM�3 zM#��m�.�
9� ���(ٗ.;���JTv���H����o�γ�ha��o���H�RtV�^��B��ɛ��*N
�ƍ2���l�f���Ն gWVbT+����р_Gf���D�ݪ���Ș&����Yk����N#!�ι�IjXT7�ʅ���hxeaZt�ٲ��~W!�`�(i3�?�JY�)�Y`��jD4�ݚ�Н�H�o�T:}��d��-��!Qb�Cɪ���������-����!�`�(i3D�wP�/�w��jJ�+�rs�i��]S���D�'�)�Բc�<πV��;�¬pX��g��U-�e�(}y��YmҐ�̓=�^݊1�m+�D8
�:qEp'{w#/ B!�`�(i3@ E���߼WaU�?2����W��_��	h����QR�^Ƒ�Ӎ��t,���~��;�,!�`�(i3���F��O��ݚ�Н����F��O��;b�-�2��;�P�t�5W?�;�끣�os�鮊F�7������;_��8W�w��fD���5�Pֹo��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc"��`V��b�˸eT�^�KGUrKp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hS�r�F��
�@	*�F.��L��Vy��H��w�1T}��<+���SfE�����z3)�d:5�O�%E#PD���D��Sw��h��5-�`��8�4!�`�(i3<�6�Q=)FŒ�J7��仂���Ȉv=�¥dٴ�]�!���3��L�F*D@��jv��9��H�fі��b!��u��	O!S�E�q���U�!�`�(i3���y��lD2�û����b�N���޾��(����T�G���,ͻ�������n9���)��=������c�Y�{'%s:3���5C�ݪ���CyW�f�tГ����Ѿk��M�!�`�(i3!�`�(i3!�`�(i3!�`�(i3qJ;���K{c�8� �.�4�F���4L"���Ǟ��Q�)F(���o�`���;��|B	|_�/W����ݺ��Zj�-%f_��m����ϏQ-+��B�G!������K���f�(}y��YmҐ��;�¬pX��+�_0c ���m=��}q�3�\��φ��<�6�@a� ���N���cp6Dq��;���EWr�(MXdv�d�٣���,�JL���ƍ2���l�{y����i�q,?5q�w��.NG�*��6��|#HK��A(�c���_G��Hb�8�u?��I!�`�(i3}�gv�oE�[��s�A>�xw'��M�v�����FK��|�H��4"?V��j�c�/���q���C�3rEe��0�U+�qbp@�!�`�(i3g�"��Mi��(�����!���|e"*qA����6\�4�@�� �-jېI�q�������?B��#Ɵe�*|�÷�Wе !�`�(i3L�J)���� \L�1tSjv��T}|�[=b�͢�7�H�Z�cL�7�ݚ�Н�V/loo4#Fػ�ܢ���|e"�SENan&��u�Y�KG�S
��n@V�� �9��1�Z���=���؊�9ب�ݚ�Н� ��ս��	�|�O��(MXdv��2���q2ǅ�|0<!�`�(i3fF�5.]����C�i��^!�`�(i3�ʃGמ�1F#�֞q�ƕ���f���fa��zJ�r��h����Ơpە|����<�ʅ���h�&�(���D� h�ҩ��wӨj]h���)��=�p؛'Ǵ�'���Xw�j�7���W�6?���O��R�^Ƒ����"X��[��	d=�4E���b=R�^Ƒ��_uc�!�`�(i3��jVѭ@!�`�(i3D�wP�/�w<eп}���=��Y�$��L%�G�b��6��	㎾��;|�5�%]���U����z~���D)9W !�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��j���p�@ 8G��5�K�b�]�{k�h�+�c����`�1��W[ �['�t����L2�y�d/t5yz�N���}I�^$D���p�n��|싉���1�Z���=�"j���b7�m�e#e>�'�V�k5j��Lc�u�f퀔�����x/<���0M�����������@�a��
V	�){QV�*)�am6�B�M�5�,�*�ɉ�|9��r�#�SfE�������E[ȟ}��ɣ>o·,��8jӟx�`�G�v2�\n�=G=kGn��C��k\����K�����3(:�QuK��E��^��\�=�#Sh�?ҽ�8ᅹ��1ϛ�8P�tK��+�(�QE���F�ޖsJ��� $n�v�������m���5�7
n����F$��_�>�{��q�@�в���;�{���𱍞3ƥB��K��3&%��^[Z��E��3?�d���&�A.��+�W�QԦDN�Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�z�C�f��H����������@�o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc嫙��G�-:�N�Ò�&���m��y��(<����t�urg�2RX� 
�N���2�t'�0a�i����i�d�٣���$u$Yo�K!�`�(i3��������Ǌ�r+��M�r��(bv����>��Lqm�����*s�}F'�n`5�fK�3L��'9!�`�(i3�� л�������@bpVXR�CpE��:���~���Q�W�����a�ү�`���;��|B>)p��I�K�ϵQ�VKp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�v�d���}�P_FV{Q5h�nF�2��D�pc�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�$k)8��>���l�����G���5�%]���U����z~�����~�r7��Hh�WaU�?2��E���b=R�^Ƒ�ӧP?��;��'�F��sߙ����pz���t�T��?E-h��$^(?��"��K��N}�m��{���q0�/)ONcx�:2QYeƈ)P<�ܓ�YO.C�U��B��-����REJ���}����Yk���'ž1�|�'����z.��W��!�`�(i3��4h�=Iz~r��V�n��dK�����fF0���2��}��D�o�&x����E2b�z'hۉ)��d�7�qĹ߆�p�h��d��JXl'�T��~��?u��C@<�6�Q=��ž�Ć�T���7X���c�}��
�t��T&��ۥ`�M?��y�!�`�(i3��t#�V�g�Tԝ��}Dq�f�5�����}Y��	}�@���	d=�4E���b=R�^Ƒ��QvN0sj��!�`�(i3��B����U��n�n��)@�])�#����9!�w(�y?
�:qEpCt�w#��@�����!�`�(i30ȉ?��b~*��sং<�ӛD��q%S���Hd i�rj�I/��\]� h�ҩ��wӨj]h�7M	�\���!���c�A�L'0#P�O�Z�d-�~EL%�G�b��6��	㎾��;|�5�%]���U����z~��7��:��}Dq�f��	��x��ݚ�Н�?V��j�c@~~K	�=��Y�$��L%�G�b��6��	㎾��;|�5�%]���U����z~�v��!�K2���aR�!�`�(i3��Ě�����}Dq�f���Ě���fR��}���;�P�t�5W?�;��׏����rKR����a��~v�VV��	��yݽ��VR�!u$
 Tpl�o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�6<���Y&O�Eb�1[��?��SH�6���b�O��]��Y�g~[�#�X���ħV^��.�v��7mTp$���"����\;�e�k�j�������Ky����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���X`
��Zi�����m̤/\�A��������	(ݖ��Mb,�||����~ q��j�J^2Y��kک����n|�p[Y���"���E��g����X�S�
nЯ�O�!�`�(i3+Ώ1;��5�}�]���LVm��8�`*��*!�`�(i3��?��%��h�r�Bi�v�V�f��?��W�
nЯ�O�!�`�(i3+Ώ1;��5�}�]���LVm��M�]%�����X� 2!�`�(i3���8�8e[m��! ���ÙK��<���
nЯ�O�!�`�(i3+Ώ1;��5�}�]���&�G"�2���k4��X� 2!�`�(i3���8�8e[m��PC-��i0Q�͹�Ɩ,�.�&�8-�!�`�(i3F��|�'�&퇖+rv�a�L����Z�]qDѸ�3���L�l���̫��guk��� 	-�	��[oX�;�q"�ư�6��lY����;AD�,#��N�o��f.�o�.�3�O�^M��`���O�DXt�ny�B���v�����_�_Q�͹�Ɩ,�&�S����A�
����!��Wݴqz����H9��p#�7�4�8Z����